-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
poJ0NkZiPXNTqYzn5erJdbx8jxhQizsWkc/6e0qnEy3agtdQM416Ggpc7LFRn3RevKA64Qm4ugAG
/+tTeUGMeZ/Wrnc1WzZxGrtUDLImPngUDnJSIILGIfDOqSezrYvXzMI62Nn6BB8Qh2fguTM2EEh9
J6dok1ecG41qyVZmCeurXCfcBOP9uZlbJH23+NlKylLjnMtsxTGLRskNg7MjY17HNDv5MAL60k7T
Qu/BYaAh7EAOMW81e9rf4BJc63crp/7BLqemqa1KnohMqDIbipkTOV6uOSArtCCKxcrUXw5wQ6XP
1GEk4pT4eovTr9qdfD3lvDEOrhAlxmqMyOBt4A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 11888)
`protect data_block
6LynMkTja5zKj3fO4IyOqdLB2jqyoGaZFSlxW4SdHam6/qbpDsAP4o46TMYogY0UspkF9Tb7u7Bd
n8+lkDldxCJMbS2n5M3oNwyZbUf+13ILO75y/qr0ZDjTpmReIVSq4MU0vc8HZZHLVeCLKhuHH6wv
+5/uu/gIukKA9dWeDy4LY97QMeJ74YL5QEtO8vWrEp52SwNEkYQ684LPXC4jLWxuFvJpHLvysFpN
gxDI3NIDWVkdiSxXN3E6In/FZrQYu0sTOhsvAyHw9hlh4ZooBjO0nTF/htyK7cGE6/ekACXEiB4a
V/EF7edNDU/pK4vzDHmfOUGrFcQFBwju1BZQLtZfo1NaxTHSrkE7cxl0hFWZzVI68ysx577OhkKs
8My8ghQIDaG9EmlUUFnyEKlIaru6F+BvdXJJqZuDqr62s/fnzbBpLiBhtXe8B/9ZixEfmtv+UL5K
9zhbRGA/w0HUb9iiCuOUCphwUjuaRAM8VpssUiiYb23S30dDkEB8H3TQQMRTH4I0qP9KChOszMLB
Hc21t5q1U0gZRVVpoaAq8buNgimQXzjkt7/hopMglPtVNv7symvUdVhZvNOpvHJnhxrPOq6ALf2/
EEs6EGJbgPkg3ye64tBgJC/NJSEJsQ1HPyXc/0IK9ID2W2oz4fnIaTJxcD96+vXtnJHAESSWGeI0
pMYcVYmgK2PymEqxmnNMeTAD55RE3LSdxYcQJDd4zevHjnjAGBssjJgoHzvuH7XUheM4nH9S/rnN
iySW7P5CvQo7mst95l4Ktd+MVnHXB9I28OQIepXQEhwNGRtroNkdvArewbmeKAffWrdIr4OXSsht
RydRIy7ZtjxwXXi1BokDZoYJvJ7OhC7xQCgjrJ9pJ+gVIjpRIk/+0sxrh88qklcjZScvwGtgz95V
vn0Pad/vHye11pz6GQHV7jCJaPD59Q+t5Mx32VGeGTmtr0GqnH/w9hehXwW/f4koyhy+tqWCtgF5
rP+sekR0GhMx2Zjy+A5BW1nq8vwGXgHSX8M81x12KZv/PexjEFSKD4T6eUmTNvOapqauNIbI/vJp
6RzGxQEuTYD30GGRpzfcm7pOx3E23/5Sg2JGbkXwwgvaPJHbb1GivDWQT0hYT3uNfeIo2+/G+7eT
yrGzrexS1/1t6n0XlGRCOpyWOR4byordEarLTX2Urn1IL0mWMFQK4vFGS/BdAw3TVQ1Wca3PVYNn
EiNAlCtar0LWT0TPP2RHSsbVk8as9/MCvW9vFx/Mrfa872G+uu1YlW2nDnIdk6jUd3U/2UL+qag6
XJACVlLi4SoTRwhLeHu0A7+XczmZHSTAHRp1QzHPBy/r36/IOglYl5w4twSp23tP2zRPgLRtfTLq
maBXoT/rR0gN7Fm7ye9QTZyF3X36vwwl0DR2/XDyHa/9ta1U+Kb+JqzyOJRq5hb7O+G+A4tIjKFX
gZenzCxARB8IxaaxnOs/SrEtlZraJ6T1alOJOKfls9vOafPVFqnGGk+51FUCIGg5Sv4BCA9TpZtD
fbmB8pOyIqkdgVGUw48WWDZnXr43s2fvFmFNH2VHHiCXMgYjboLU4IPrkf02eSL0qq3T6hyWoyIz
puv6SnMJN327bsh8bQ6jdwWKHTwQ6cWjUT97KJAC9mnOAts0hRO3kSXOtVNvpL+Z1Z/8eqvhf47M
ztbUFmI8qaFBi2SNf9CuK4VGatMxlKpXL2ah92uXX1KiGqjgO3lQbKBYPj8uAwkIqiUJHAcse7t9
6JaCRmw8eatfpvRW1tNeVTdd8dVkRLaKRJl0fyZArYxpxFh9efxO6YGj6g7KJIPVcEEf4Vt8DO02
BgdjDItEhUF/RUPcVZBe+GLJPigBn7LyrYfy65nBo3vQjMEfjkOqRmj0wXAifNKVmzp+bkA4OfLs
LEDFahkECURquIwu3D8COZ1Dz9mEMg6YG4Ijb1d4r26r04OSyht9TX38I0j+tosLSozFAib3p8Uu
768YYyZRBtzW4ndLE411tjnYpHPPRnTPc4qK4gNO+XKNkLseDWpd16sgczwOuEwTwyQNlEksUU10
0IuKcVJnidHL3x3BnebiYSKSARZrdFOxpof0TWfI/Y+ZtG7RzKG6IoCDaCNdnwAejTLkFWMOvjMc
g2JSNV/a7aY4dPwGlYqFssULoRBzIOPjj2WjXffsSvnxJmEvFDYsln42kf85e7mtvL6eR3bIeAeb
wR0wCuwS9CD3omvCCDMh9T6HqnZ6PGGObWXL7tGga19/3RnBMpSkV22o5UEiHH11n4Ilnx+gXsvA
cjoCos+pMzJ+5k3mGMp1HdXcXKSPNg7P/cxC4Vpn/s8/3mi3zc63WvxdoB3l6RVZGcNG8Q4rgdiw
+lEF3bFQhyahmQW3h2M/H0R1UO1dLl+Wez3giiX68PP7IQKvW9kTbjemLG1gnRk0NF0wQ3cj0161
5/WvAKKTIcqQdBSrkKZKVZ6EGv3fVE4wZNQ0qbjIuhWJSlRD/vAQBLoFDHR20v1RQXIgNGSi8nnI
MsxerMSoUPe+oZ2InvEeh+4lOxl7kWMXnOuosst0kp1DqhnsBSiHX3x3sTdOSyoCViy+gx8BteAy
ptspN0iNhvDVJ4deRiNFzXLMu/Ntm3V5sKA9rNUcxpcsYcCYMoG6y5nvNRcN21JOCYV1NBEWFzoL
JT2UaOGFsU7/oliC2f/EpCXWTRkDYY+JNkTp01AoOglzstEsxN11CqHpUBwARs8P3X4k6lECGW4v
xhVeIScJKS2PhgAweo+F71YtgUTcaq1Mr0q+zegaWAXpZgZWoRm6AvnBGLwqbdkGMMxK1GSVMlCi
kvXat3m4IYmiz1zIs+27v3UEgNQ9K3uzWVcoTmCTgcNwzrrQzYUhw+glomktp2tFJpEhtPW1BPRD
f6D224IZnmUUVVWhcU2hT6EfUfjaJ8Bur0ceZ8A111O7YeRZFEEzWMywUq8z8+hLpgz2T/J3kWnD
7MwEj5Yr3n4kE5wdAGoIWtsaPZ2L2l/H3DIw6HdARxLZSK3gfCE1yO0/b4TS4ClPhlmn6sEeptFR
wIiUaoStjkkjhpRxgGJUHF4eTeiBUAPvOu6/AJ/L52QjbLg182mHSqwo2PNQk4v6z9ulfHQvmQbc
XgyKPVPJIIhCzaj2TLi1CvNHMJ0X+J2HdUBumEFkvmLzRfrQDnfzArTXC27TgFX8OfjmJxTDPJpe
/l4wqo3CSacMCzqd/wLhRn3pjFTe0WY1k4pu+4w6b1LeRHfupFiwLiGYgr8x9bjEaUuOIrqXClUA
pIXctUX7OLKJtg5piFK2F4ao0qyiu+vxqvN5NGQ27RK54JmozjHDwfzZNlrijUzLpjm6S9lRqDpu
Xx7l2l1xCqaMc91YcV7EVAxbO8rIHz9NpuUIAv/iwmlICJdfLLIsBLVgLRabLvQ3iO+JOYmWv2mg
vQNk6b/QK0L5dYcZvCQPCm4qwvDX+kLh6m+GJfhNXsPcRpRpmLEyaCSf3EatbyHH6KqorIFmfi67
EHAEwQBg2e+3iYV1Axlhotzmyv3w5t2P1gooy6GgclNF6pVnC7yMQC/Fr91ONq/Qyh1tPwpF6q10
0jasa+HjwoHJJfW6PjCwN7RrmFSf8b8wkeHKM2TBAqvkEfwEH3OrEG3YjVbygLcr5tSp3b5T6yPG
7wk/xXvVMpNx3dz+r8dG/ioIf/xBYW/c5QIKjqIwt2Gdd5Zjj0bgP+ymCc2p14BmOd5BbeTI2MdK
Dnt62ZDZ1/KuDEkvuT7iRe2Dem6dhT0vKzHu3NOGZpdRCAL/qs3WxEa9DuwXeFO1AYnQoHU+e7jC
O/rjiYnHID2iwMW/rKwvI60zDf3caj9WvljcAUzbobdygJU5gR7IJE9H1V10/kDsV4IhfKrjK48x
7TP6s5WHzeZK+5uVhiGt1PWstcgPUKVtEWtSUOw0+dvlTjg+zxnSPjB/c6b1nIERUkiAwd9ysH2k
eOVo9ZQXqoPuwPqDAJMF4tqcVXPI4Fq81a9LsfEIR27PYVjeke2fkfH6nMwqwPlsiWkSS+YbYVMS
Y31Xhn8VQt5PQV1HeHE0tGlp95c56L9/H2wpyVVobr0j4sIzowd2Qf3+eGK6bwifHRAPaMCOvsRm
4FFYV9jJcydWDD80Tj3N46n4sw8pfvEyGOBW/+jn4Uq26OBXBiosEyc7r5qD8ywLN/U6reSg6o7K
y0sEFajaE4czHBi5dh9hebzUrhq41HspXy/l5xl2Z8Xn5C1JpeYpAar9uSXaiSTtNJgkSUBTzw9c
ZUVljhZiS0jPhY/v75vc0KVgOvvQq6ihAH/Rnx01X/OgwICrVOMPKbmOgGmJs8+PavuzZjIucVxI
5gVPFfUtftTViIbVnoCwoZT2DreW+V27j6ZUprhtPa+Ogpwpqbt/Ak0zu/oVK2a/JlYkACId1d8b
PUZlB0zdM2rB/XnaJRaRSfmgC7SOjfjXAfaHVcWieYvMF89mqN8BHBieuFsqcKFo1r7oxfRipcqW
i91xma8Ag2xrCmaoxZ22cdL796h3bJaGKeAuBVhgvgMRoYfr4INYl5Em9MA/pz7ELOyJL61OPGbY
HDyBK/7p45dEM5PDwbOZXLS/JSYFcWTAYCjapUc4vSv8eAFPwVbkTNSHI4nycZ0wp8dva8qPMTFF
u4poU55sbrdfHqV+E4OxaM94C9KOmVrwCnIGsoyZi6NwYQc07uYIhOk8uYl9FYpfMvWJTFZMMLKD
vYDebDwHZq+rzJkboWmCbZbgr9xSFsZrzDtIIdevMu9W1qZwYgszSd3gRE/SG9uj6rNu1Wbmo8ol
BC/Ck6rxVGZgrC8sqpM6OwJOzmiHuP/HOvLmVp02oWMWu5XkXbk+jmXKMb12o5Doa9k8bR8SrQt0
gVDVKJOT8KCzwJkyqLbVsgRncGQdHEWtxgYl/8PwMSLenVKgjFhtwlbhSPBLsAB5kVHAjRYdCPPk
oWwH2t4idZ67OvseIUITRxnym1LLyXOa+oLVCFuxqEeh5NpWtvkrsQg40qF4uoFpNFaTktn3O+dd
NIqQTR8RUTnnya7wQBMQ+9Pwwtng5bRoVD6hUv8TbnFvcY+QfcK8n5ZRL+OsfELyE2Pp0LuD49Km
6dDBMeoggy73I0lMAYFuuilOGOZDa/uV7jBWjVlwwpnQ9ijGaOlpOVhrzm5wlWHHZ8P+lW6bKMhL
WbtM7eViVs1+AgnM5b7Q5AAtKR/QA6uucsMS7M8bklLexjW3fgbx56LWb/Cgjjvzrf9eRjbfV1iz
mMMC2hCcqjnPB5vdt8P/8ABY4Q5PuroagIABB5SzimRsWwm3nAdpxvGs42idZF1l2ZBFVJTJv6M5
1opfhZGJ33xBseNDbKzYT4bIXFyFst3UOa+Q3lsOEVGr1U7YeeHiYnM9Xd7VM44wtfahFzmoUF4P
Mb1oyl+aBKQMwgG7+ijgLHgBXLRiEpDo3VzzQ1lGEJEthg5nnGMFwp9GT5lfBFYWzqN2mMRq/Sll
hGErcdZTcm21AK1HpC7RxrnYXGxi4BrfX3WURBZ507RHcyw5ndJqMm2TzR2flpJvsBUZ5/8pugJd
e3f9nUmtzwLWLq099lgTYtdGEwFxesMpodQWvXFREGDz8Zyi9HFnBUX7fL59MgyANezaUSXGQj/c
OGBfWg/vXA1C+9l9koYoECrv6NP5LGQRRWgzAA/1Lny/+KS4GcbeGt3MQzHa770PjZCJy0UEJFR0
B3/ZH+FXQfmfNfzSIglpQcM8GCFbLC/j5gSRlyU1QXwFvmTcdzjnbIYPWQp8RVyzdZeC9Jy3DZrL
BEN+VtUWk1kZgaplSk9Z0f/J1Wk4Si7yGu7uV5bPTEyo0Mnwn4yhGrfMmgh4to72LYTutNoNK2eD
vo5FW2m+x2nxDlX/snDDPF097MvYOWXZ9evTxXm2iG0dXnqHF69NkPs/vuc1J/RfltRy5EF5Iwh4
QsI3VnueaH5om1nIyLsRb5jJmh7dHE6EkNB3en40MkcmbLt4TXAXqSzZwXkNGgbSssWgS3Mkz02A
gY30EwvC05zvZ2+R3zNbb5VPm4+Y3VcI0FpXJR5mbjSBD5hwwqAwAzogDdVIc4TBySPeXSpTccOP
N4MT5k/+oLWLf+0g5ELvyc4Mvuw2dZ0+L3xHfF0yR86AdtzgVPiDuY+zm/lAyrWUCQF4CGBDytvG
Zs9iqP8iCEUEuCk3Ib/b9c8ghvKQyK4Apj+vNy7b27F1ocTK4Lyq+NXdb4af7AReWAFKZRpEKQOI
L/U1h0Pm19oRgJPMB1SKXi5jAqXwZoQK7+fwRxg/0qv0u3BmucfqRQkNxsllXEJofLZ5cSiY1gmJ
v9HjvYi72MZXRtfwkaxRnUoJVkVCYnxnlXCOXks5+kxUvPBbolxgXrqrbG9KMmkx54AK/1h+IB7d
zELW8K/fw/jDa7MXV+DiJxGklZGVDRzlO+a5G2nvlGq7R4F7jUPIlSbQfkrccFAs2LPxhaJZo84x
UVXOClTRoO55VjSklmM8O4bnxtjY0/Y3TTSHjO159xV/BJzE+tX7tO3mmssKXnxsIKD5CP04YHYq
e7Fzc2Ob6tv4Odfv+M44cBGw2GYMzJ6Z7IM5tuqDJvUn9Kk7sz2tRnEU8wbgUOE6acLOzFrlJnFC
9yekJzSS6xQ7p1wfE3Jp4KjHEBXj8shS2a5o6GWzDHCfptKZhRIkgTRA1PXdC4hIk8dwYpjtC2/F
r4qbBWQUKxzMUXKUY8Bt5yWZWn645vjfLPnSJn23B3AUJ0rQb46NjhPEtehrktlQScio9zNg62R1
sJldmiG4oTE1d6zBBqJ4GL2/QNiV5A9YPCdnHXoGkW/AM07nqFuf9WSrbCMfgyLAWEPpSs//7rFV
wvdy0q0HZntoKvJkLEHD2L4h77KThwzno07Y3ABMmI5Ka/Hj/+1xG4K32PzfyiKThH4dgrYd33eG
nBgCqdGg2fR350Zhw/BLz2RyYZG0S0x/eVs+VXjN5MyTOyjJ5R7d3keimMu+F0Lw6ztg50QCMmVb
tzO6C2uho/qvTccgxe1zciswCrbuqqboWHvm4tKIIhC7ccsfmpxMdh5j8Z4IzgeOcBhpiF9MzaXe
yTtojKXa99nybcKlyRIaArLHxi9qRd2OA9vE5qJr1FE46SnALNUFH5frXKXmh6HszQ5H07xJ18+D
Q1ta+szWitu9R3fj4WXPtqvRrvqPHBvByNE0AVkmTIIHN1OgtNSesfckUixzWCKmJtjrP9Uj4IbI
w/qufSMhIKRnnjdse1W/y+KmQ5qAjE+tF+IgOQAGAiT1ICanvQtKKrVRb4N1oXTLNPrDc8K3GLeD
aKBFeFx9fcBJQIOFo4qs0bKhLcOMcZg7fuzO+XgQg9s2qie8v/FqiaGAepe4rc8GOgg4NdnH6kte
elcIgaq6GQFhQQvQiZYmPoSKvI490Q5Cpcj26cOwIPtKCZw2X8gR/zF8Tm7eCUeszYHLBEYxKI++
3GRgLrIpYu8FfFaHKnON7DjgJmYcet6VkXeonFfJUzIYGIsFBC6/OO3uP1pBA1yG/8oZGceBIE0z
Dj017p29jsSmmEX/14Je+dguFq3WvrsLyzqr3Jhz/PI7x0J4f1PFWlFHfu4tAFJrHX1kWUi1Mdoi
Cwuow2m/v4bLQl0ietqbv2W/MwDZLsdWd46VTSnvVeDJDS3PhA11U4Ypd8E/sHleyVv3svsGjFCn
8q4dy6nO3GrTKHIG0V4Rq0jPGsOtUsC7kWS6GWQw0aiTttkzmQp0q9T9e9DfACKDxAezADKsKV0a
m1MOcm1yoZVs9rBzk+marcuJcpXYDOX0Qwa0Lux2fN/smky5vm/YjqPKNUljgCVghHhSYuTZ4dKa
7t1M7dSrFNDc4QiX/z1QCW+kg7Y0/j3nylHhj1f7QAqflqOWphJGjdFKaKjoSmOMzzU/yyEXoVXi
+guEAQ15Jl270PQk6rMly7ZVxGjlw+JO9/pPK5XCyoP+RdW1Ax51MUWjkF0vL1tfx/0z3LHGDHUh
rZR5lk/IgZuSgKtWTY8JDGEDak6pMYp7xufPDw4B+OzFOO7BtsKLxrDnRqpPCdzeFjvrWPp5PbAC
bEl3Qo2V0Kap+LGYKyAJNS2FUXYPcYujUg02BV/G23fFJx7BpJtY2Gi6tJeELXsL/ApGqg50CNQg
hMXqegVECjySz3SErKYTAm2zoIXvKqig/R0qjeGIGqcFL66T+/utnltsnO123/waLgeQws5S9qND
6c/VAubb0nisvtDKJHqWKqZOMNgUUy0wC3DTznOHBdSxNm4Rj7H9DuAEH2ul/kwxpwf2PHslM8jR
BX+kpvv+KNarkIsYTZxVaQxdiwUULvHQ1yEPijTWWF2JkqGFDxFawAQq5aZ933+Z2CIBfrm3ikTn
rSQ0lm8QF1XlhHMZiYCHsrDs0ouiNmqRR9I2/pb+TCpz/RWk37THAYJj1fP9lqDxT0OGcwQxrANG
NdvZhb3vWVmw9ziejXdTqfZKUnTJlUF/jz1Yx8kvkRXWaHrDhMtdq92XwSaAacidRhhURe/NPIsn
9+V+VFPVXSIiG7+MA3k4DVMyJDqZhJoJxBZkOkaChk5aH9AcYDtQM3Iyz9ALyrLpror7dlpsPJY0
rOq6js6mmj6dSct5IZ3+VMD2deN2ZT1HWbZZfpzTwD+1FH1sL1ZoSi52B2tdB2gwD634oKKIkV9s
CpjvyCwKvSt5w/5OriJObne0laUvC08dlUbOEhHwpIMnMn2GoxjbawcO9MoG+2lQlu/Aglvj0va/
mrGizrbMguU7ZrlnGCcvOkLH+9cK3IGDKwu6AKpN89G/fKg70Qf011fU7uOacOXifc9JF07V8HlR
wBkL6kQvnX1lIsrJ6ci1/3J4gB9UBgRBpvZzWZtmeKrqB/SXS3k+5VcUFecrx93G+ClL7le9Le08
fTRp86QOt4RKg7/oELPAWz6lmNULM7CUIJs72IqT8cZEx8dPc/+9315F82VwyXWLqi6EiNNbjU5W
y86DQM82rOHCnOiXKqPnjjCs92E74i9Bp/ctp7tUYE2sLxCcenQmsQCR/gIoAQ+FWhSnRbIpxcRG
Ykpw1EatKXLsk3EaXKse0PnDWgKm6Fzg2bPpbHsYqPrF8xdOXIBxDub+yU9RRhf/8UAV/yRNlVlq
a1JchXbFR47YKHPbN8FJeThuKcAaIab5+KykLETKHYLhfZfjNbZYeY6mfj7wR9oF/8FpqgnK8Su6
yl+dwMP1yh4iQOwKv63mgb1dBFZ8sj7uufW+4zNTtFwlUNoYYo8IYtXScmDRQhUeu/28Sa15BmFZ
m8xI6+y0b7oQOtojwzz0+2DMCQBGjI5YsK4EdT3ToCAMmnng1ONArxAIFf2t8c0p4t6fPKX6KJ6Y
PNn1cfMvdT9N9spxT7w+ali58zovnS0WiI8bZ1Al/rpQdamYJILQ3l2RelEgRg6ElaLTXl9EtR79
wntJ3eyiC/o6EOx684dE4CwLnfpCbJPYZfOL7TxtrCdvscitCl7bWqGQaVRwMDanZeiv1gm7eelJ
EnP4zk3Kk0IKlweXB/Z29YXlP7kWrHaWu0syN1pSCkTa6nlXlef0adk9P39jL/KDi1sxO8fe+tVy
iOvBQQ6VcBSzwrfkI+gdOs2mVEfsKhBZcHFVZUg+NXpb4EKO1A/tvskD8d3TVLPLBBdt9s7dte03
68lnDHxG7g2YOnDFELxOImIkXPuWl6e5UWLZ5KYwCdcEFZT4WyVVpbjJJw8ml6oA0v2pIizib5HK
ixggjcTfV7SzxgvbS/Rh5Dlopq3sjJ32AmVZmimCjJ6Hlps9RashQ+LN3YWvZgDPNVI5v936FFLw
HCZK9TReprry8U5oYJO8eYBKt2ZOy1K3aBCtAC3+ZhpMjIN7VJxZNYgepQTibe5qD7D0SuUW1Ano
8KLzntmdWqkWio38VXx6ODGhBqeQypTKrTY+0NonZjad/Cu95zE34xNwC9dE2iZglwCn8Xb440a+
WbjNlBfDkASHrVNwIveqfHmspwN0kYAmcTpsa7SNpGkxWOgHes/eSO5haLPC6Hc1jxqQ3dpFmurF
eWV00OWsji7o5MVdhzhlxbIrVavFBwZRSG5MNXarEfpCKGUg8fwgIVi6jA5I75sigZg3Ft+Xs5in
vuSLKo9ttcVNRzv1t8IxCfN3VjM2vSaq97Que66xmkU0VoHsll7EYwr0OL4IZCGJBxfJ2MGEtgg1
g0ABUICUonRLLJ/52GWEGX6YYYR+NU91Ac4bCwFBtrZtE+xk4EKduHG5EklqNSYKuKRlDmjSaWak
zexOzaZTeUh8io+edLC0aLIxm1otznOxoi6SOMa4IKHcPRMFVNKvgUq1rswzgfLOtndNzTThweaO
EC8+RmQJMXqXu5G/+LyXwi6+XjAEENfFvL1HddcjBA6vu2YPY/JOps+3lx9msNolN+qEXFSTdt8R
6tcFRetXsoxGynZ/ZBbgNIRaRO+Fmd/P1qeq59rw23gL+sbJ96Vs+oNF8Uz4fCTbnzWXeTqQmsO6
JLFjV8bMwvPhstmwaC4cuwP/OamlRUY6MdC68ZDBOkHIXZalCqYPecqAjzkB9HJjM9JzdsRQ1O4z
weiaMNOEVSPIvr+utfM2Nl/r3Bpt0rfm+3rrj8h7JimRq2GFIs7T7bG3XtoGNMDSd8u2GVQoXV66
2ExEgrOatcmODVSPQdjQIj9pbT+JEbiMG/Voto0oVRYUmz+GnjIqBw9nWtQ8lJFSpHkZnYLkhgJJ
HA76KmAqlea2NidSwnGxOihXfnb1B9uZCphkhiOc/fMNx92odkJfsuNHykgMJQQ+/PWCUPUCi0nh
Grtf2g7JZQOu5sl+/42XTDqPVMe8gVLs3OeW/TvxXYkVpBdyyKrGj4jv1qFHu/SfaAtSjo+7qKmU
3fytRDpMZDZ8rXwiEc8K++lLp6PzDBMyUHIoY6nQAdrWxIc2G3ehBDQ1GsPg2kBbNHkyfKQxixtN
+9kvDPGqPXagpw4P/9bNbSP7mS2g/d+FVjgvNmWi/xP2YUfm5HyqWEA5QxBxBxkIsz5I924iVvpT
FdUVdmd0KvHlMOpPxzAYbkPRBibRSOAB/A4TkBGQi19XuJUuAYdkZ5DY9vSl6RF/4o3YwSGnFlxZ
85si3XnSSa1vLkMswpjScKzeMfKsZL+sbua43RvHVcUzzznjhiRsxxwIu05+438HjUIxHuYtjmsL
z7OOcvtBbQML+8YjrCybaG7kMHS8KeX6InYd7C5bkEopPQm6PI5hqS45avBX6eAC6oF/Lj+94TUx
MpkEah/Am2EC1oRq0SCeNQurCEptszYFAjCae6cGtKJe0CgfdzWA+TQIiDlzNUIeJndWX5Xh8MZZ
H0OVD8cpOR5ddjZfICskAj3AmGYKnSaORsab79z4LIL1zhx0HYo6hNpKxzCD6R0Gfn6cjRehXBqF
LUe7r0rirlD9R0Gio4NMyWgKN0enY53XUvgTb5eanIPJzSNVuAVHT96Rnlt5NTAvfagnwi0VUzFN
zorMZ8sbIMLy3wD6El3ats+fQTE8fv0HgJOYLctbDvXDqRXhjfn4qwUz72IqddHt665c1BDkD1Ns
kaZeckSHC2sykF21F+XCtJ1u8bBy9bOtpy2vtVnmWLZLu3hzk0bjAHuNLD3w7YTFL8+GYE1rTuNS
oqzYVGFOJSYo3+umtj5Hx+RATBjoasxn1g3gviUuyZy256duJ1nRJ2+OLq9Vakm22n3AGQcgiabo
0OdpM4P/7E3E7g/adPn+XOhTCM6Rui5ZHtqPwmaQM5s6rD29C3ZeZXihk0vDUmUYD9arScuDrcdS
gspbwOiycHWmeklU8NsWDG3FLXMO0RxojqPtHsh9r8ysQEY3nxIhU71CovNX9Amtpj749h8dYKb+
It4gWpil7VUQHfpttOqpOu533RJ7Ft+gQkzZAD66zLwyBf7Yaxhd2nAvLf6DAsFL30vSLZzQI0ra
w2A/yvO2/WAEpFVBiYFrN+lz8Xg1q36pw+eRFKvtss+zCOAHZ7EgOJYjrWLmVWfcUNIdTSENRdTH
rWj8wmN2MPLNnSKVVSEdXQwP7SPNCWjYsbHGqMfLA+uIucF8nHe4zfIz6FrBQX1UiV2+Vf8i5JlM
jJMrhmGZeKo3SI5NQULKu4Cx64Fqi3cp7LQx8WdIz0owDp7Y6pwpKG0MP+MVy50j70yyQtAP65Ce
fhvUb9oa1id8vpJ4hy3aFN52FtNDG6UCB6fKsl166le9cX0XKp2neztvFEZ8h2kIQkhuJzmPP0+1
j6deuW1HtEmCYCI3rqT6qLg+OOjDwA0xw0lMlvcC1m5vUWFP7tQyxHogLiFqObvPllCc9ruEAZ/6
EbqtZTi/gstZnsmTMl3kIWOXMYzqcQsq3FO4dI7bEBqzlRPGoiGrP/IR251a1Etzqyi8ARfC2NXJ
Ax47/s04i3cIHrWNVlPZZhZ0/9uD6L758Dh5zb5Ee4KV7xiOJNQrh99ZC0NpZ9tO6fKwd4Z1KPvH
qlDXDbipS+5FWN+PcI2TbxPmnk416JWbYwd8vh1lldgIqgoPYduzhk7mFMMFsmtRRg7OzdPfuw6k
XTmNV1/6QI3fQsHt82dxOH0ClMWYvWnChaXXxx99rKOxgmmRLcRpH33euvXBC3Pmp+E83rmaqjpz
RfOq+mZ3Y/o0S5sMBXvpdH26s8ReUNDsvtIby6QkUAll5VtClwzHYhjh2232cAEHnzBnQYaJwaOF
B8iImByrGjOeLJxpfzNsCL+u+ccZ7yrrkLOcqNkymvUNBRXSPn8dXcFaAJcA+Hc3vN7Sju/Eaose
9oEYXwc4V3UUaahCVL1ORFiKKhaIMMdb+DUmLQzQhuiPmCJUVo4C5KPXg5SSPwHSo4HZs2d2IbP2
ZbtFvUKDrvFjDF6qojbcqORxKX71P2yEJpnpdK+f6uyO/YPUudbww/O9FVHQLpoj26Iaiv+3Hy0L
MMAg9Ql91Oo6MFfc27ho2/T9Gh0nqmRgsJhU0a040JX4QadqumfxDsfmsDQ2VYuE6lUpbqOCkrcf
6ClOHODcT9gyj3+rMcN5E1nmqTm6Qpe7SWSMw+1ysTz6cXJ3xYEhykaFV5uOeUp6trLiweJAgkRw
YUnHDv0iMbCnUDqfTgcN/TXQWiEH46lnJWFSn5ka7+Y6UqDLXYPodk6R2j+gL2RhFsUG8jNU9llp
ZIyGSmgAiqu9H5r/GjVLEbkbjLm2HCGaEkCywceMHBEtBcQnWk/FmE7JNKJD7O1MlNdIHxvvVGPa
KvpRwU874l8gnRYU2yDWOTxE5NdOfYBOhDD1u2y8M7l64AP42fCrcHcYtEbpDD4hHhmhIlxUX97n
pJlVUktAKUtmuWMe0kfaIEuHKSacfZNBTJBeqCdCtejxxpd5bmd8bLh4pi9iM27IBRtViX1mSfE9
La+8yVC2BUeaINRmIcD+s5qKrNtgdku6SVJ3ZfzZwwruOdPVE7ZC77kteOAjPrIwOIwWD0Mz7mUV
KmxAMLil8FgfDr/H4uXG47MksoVIwUBAdfexI1Y61E8WK5sRfYeBIbLSQXV4XfG3WTOQ2g9d5A3S
V7T37PI2QIZzc/NT3KtPW/+Cb5vQTvpCFI+OL8sM/KEVWGbv31QMMpjo/O3zjErF/Iqp5Q2OI46s
O2vtgZPgSuBjU/d8ZaL+AtW/EXJZ8QzY9LgIJpNPocM4gkj+u/i5HTC7fOQz2Fk70w10b1ZzKHJC
HXLA0VjkvnWNZC5SehQaCQM0RAb1XBWSynKdyYW7BpK6O9kHy7xmroch5QBjHVdcmyFVZfIFWR/y
69izl0vpCT4clKU+Hs+/IOpVFJ2Nt0VxeCZOHBAFkke+tvEVGb0L4cy21/5RAzTN49mwYrsnn4sN
8xQnqc27MOEcZzTfFjOswaAzwH5lnDrROwEYlQlOxlQOR+2ZNX0YiXG6hbhJPKS4rbOuFAaSrix9
Gx3nCKnY5g0O5XLQn5qVLw3ombuOvBMX6p5dW4n8zoJB/IOZHLMgCqrF4nhthQ1i9yC49Sh1Qgw+
qCekmMZiw2mMcl2V5UeH/XoNrYk3H7Z05lWHV6Wi69b+XhDT2rKCB/sid7lYMTuW60SydaLHNdLR
sE3+UqqeSyyDsoDXAJ5FkDHZSnmT6gH0qGMmRfDyvE7Bdc2WnyRm5dds4R39OGhcB+aoBcYC5p6r
y97bnYg/9yx05V5fiSuS8pePOsIEk4V7TTgunWl23sBrPNieIpbVELQ6r7Hu4rT644xejwutMyAj
olJudoUbxBgC7fFjWdE9qRov4mkk9PgpkFJ3AdkxO089/tqUI7B/0yyexyhJkG34bVwQ6/0bAwwB
6d8BOy+RqwgytJq+Pm6LYvlGHKoGA71An/mAlazzccpN34+bay7XVe2uGBJ5XZRuzv2Mrn22s2gY
SN7H90q9bzXDD1bxY9Jf2sOmmgR36wVdrY+3+bcM84YMVj2Ho8/DoV2qhGfGwg2Vurq4phwJacqD
bfDqkhQiL8mRmkey5nvArjARPN4QVYlZa45tshaHjnw1xvAiV9G5c2r5G+pBRNhcIXfhClIIhvce
YYLgj+Kw40sP1HnZcy2D00uparWwe/jhTzW4kwcGXPm7E0DyWbjQIY3RPDnG88Y8vCm62eUcSAxL
HOkKcYT/blxg5aQePogW2mdZbQSs47grMv0pTe63LPXNqheQxTzPYw14K7TQ3037SCNH5zoCek15
JhHVcU8TFqMHuu5R+R707RZ3OAT0iPM9N4VfDDjKQih7M67eo9c1TBZ+02LIJTcXZa569HrT7Sy1
pUjpbIe3UU5P5tLL0R9ppgL7T6iHCqwyU75/FfkEKmv/Z6q4DsD0F+isLNjp6SNb7/H2TPJCiFb5
2oR59iTxk0eHXHJ4viShaQUsznvYrif8GXTEsBvSEEL37XhCOxo5H1w7fOiZQ8j0WnXhwWIhlBzu
2DqWX9HwL7zKoNL2AE+GDwtVvJTyct+Xr/MdvmAxHk2TGdK1kv7/PclkIpnYhZV9s0ITno/XQF47
C0SeLIZmuJ8ZSym9K+OfnK7pVttlog3jAQ1OvVVqT5ktpCRWn3yhRoHSoZIIM5fzXxZmGgKXDVq6
IrUkW7X1zt3ZFoFUfC66DdUYg4OA/qO4Sy9gBBYeSslYfoD2no9uW8BCSb0QkXTImM3QJuiQFoxZ
RV4cCtAbMOxizyfIsK5m6+6snBNK9IW4wB1EhCl+eRF96r0JLRxB6mBYO9uB4t00p2zLm3jVogBY
XPvb+du6I8FBg48wPak12X9jVFPP75nKvlqB22neHibAxSrguKQq/wlsQIDUGOvD9snajkIoCj3I
4PMQr9jXhLUhtkEjTLAOMU207zmxdA6pTw8bLMoSwg5b66cI61xHP009FTHdR0dr8V8EeFNLXLcx
E+CPZqB5L3wgkkStrsepJmEOwsefwDdaesnZ+ZUmhA+d5qyF/dN2VodaHyl4H4vhFS9NVLxnjeYN
9gi5LV15ubl9nB9RunsRCe//KtYroigeKnQ+uTuH+b1xFIc3pKu72aGGSuwO8vbL4Bmqe6HWZwF+
RIu/q1dIPVS+paTGHtW67+qgy9HNKEgvGfxLJjiBr0kvrzy8RrEhcR5Gs6tISvJB/yW/Stls6Age
1Bb3A1KzBBdxd3QUaoIFWec1D0RsN+QjEcxPcphuJvgh9Npxv/lc03mFqBd5626WyQNP7IxALF2n
2MP12Ykr+Xd874KtO8ZCCzfwG2F8lUywyHZTx+rW3VxFNntf7w2oqP6qpeDf0Cb4hB/FGAnScTjR
NfVW6Hd1vcYBS2Y5Zddbs2QLBJdIiYOCBPCJAh8tzMZ3w64++4dk1NoxjvOWFgV1TiDYDOANAC+b
hx4Hfyh8KroQlrSnFskaAFcQQwCKZ7dhmcWB7KxbfaM=
`protect end_protected
