-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
nST1dCRm2gYi9stbGD9iSt5xjC2ioFp8j3FNEAz7LqTJeLq8pB1ABsNW+aW64h9JkVYYVrcBWTBn
RUrH6yLxPT/u375HkZMugtlHNALXRAJFZvI9/Da3xiw7m0vqZV3a0m+9f8uG1NcaK6gCV5DXDcVH
MYkI4vuW8WHR8mLdwjpnH4c2euKTWgJtzz9/jtPeBsh6CMCDOkRFSNHE7RJDAhmQtDIuEFjDdRes
b7Ld4/JY+mFi8rEL4ABled73kOdnNEYXH2HRCxF5/YQX7qKgEvZaZB9mXWoIS2h5NvBOS/VHS+Vm
eqKBUO5OP0lexZ1njjdKLzQKgpmRl1JiUxS5Ow==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 1056)
`protect data_block
g+s0D2xYOxBuHAIqCyeLZ94rieOVYy6ZvkqlEHk9Encrqve2yDXYGbg5cJi5ogqKdbGasQIxhXfp
9ZkxjV9svZPXFlRssVbx5HvMWU4t2BAlJ0zQ6umEwChbPgeSIfxmQil4Pftuo7DuHJG7hcSul1d3
26a0oVwuw4JkHmqnv6PcJUjq7Pm3Etxh+gVfpZ+moxV1iDUNF5AqmlRkm6e30lgGCnOk+Pw9XFdL
PuhdT2eKtNJvDnJ3ZXup7sj0fAAmjpjJdU1PFeqjeUFZjKlTYbL4ajTUnhjLxRgkAeM70eJ1Vvfd
zxeFYabVyX/A2S0rsTmqTmPucHyiVGY5YRmJ2Eoqvi8d8DTvgHHR+QLR49o8R+Avk+1RhWHPxgyT
jLmrlKXRR9S/MV3DW5Igf9BQ/8B3D0oncOhOwoT3MC5WwVSTPIFZtQ4MH4Sg+TmOiTexnSXTvgYE
cXU8F7eetcsbknWMw7WD5cGv8TiWITsNlTd1OeMGzDt7nWD4qoMzsoYKH2vFIiZa8RyDvTn1eodB
r4NnVhfM9GMwEuCetXo4PuQbZQaEQvn50PwMWk1rtB/wOq0vKvZlT5hkDRJBAoNlb1XAEIpyemrQ
VihZIDjOrpzlbMBivsg69wLGuD9NiHIfIjV8deLfQR8t4gtBUg0PfTRNI9OlrYZ0GsZSiIztLV+C
BP1I1g0Ghb42fkDrrmTJovP8amVT3r+4yav/RemDGEC7vf6YsZssRSONqmUpfgSxuHUBYRV/nJM0
+u7LFH3gz11DRDYkeKozAnHp52Ja5jTEGLEzk9K+h2EP9SZjIlaMtVAusc2jOErS1GBboTssbR/0
IEIBb4kPC2SFQdWdPofZntsrlklnwMdogV9EpyoWV5asZPapkHoDaFiSvWLOYYd4cROTgGtU1M5D
35EkLSbhZPoqRBDxLoL8dt2ODA12SRjSwgpvILnH919UIuXt47qe1G49h0XD9ringYmKhpNbS8hu
z17Rnl1zlyvlSl9xmeWI7RhF/z/+Oh9TggeYWvfAsGcK8VaoOaBm6qqUdnBEevIHIo5bfe7jnz0q
LWDwNjVJKGrCCHvMZgC58PLObPLnlINa7bnsw4NH6oC6N3Ah0wmZcFjp4AdqAuQmUp6wtqXIc038
qazpr9jNgNc/sfGCz/qsjuX+jvR8I9IaHs//cyYHWOqm83yUADJBbjNeK0zGkBdYWw9d87TfSjyN
NlzlxakLtwTFXHV1XPE+Bg13Uk5mu4z6vSM23rHl3NmFjI5JxqGwZaHN+Uca9M78TaEP3QedEA+c
P/akD6vcgdT8VKsILdLqKBbYUYHAT/35ntheLeZyx5vHUh6q9qWQwPIHXk4u0KWLm49321V6yIkF
vJ/uS/dR0r3nK6mIlbDiyh6gPwocc9h2S79Maepp
`protect end_protected
