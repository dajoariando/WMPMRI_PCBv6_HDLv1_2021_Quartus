-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
CI8FV5C0qipADJ7eFHo+HWggIADudlRBvnaWvFNa8Lk9GOOCQwjmmpL+ZeDQNi/quzLaEn/XH9ce
J4Y6pRoDGO53Cy4+JCs4iVT+E7q0qg9SQyvvhAIhFvYc9qIxkgPwZpduryMv+M8gDKsk78W8EOfH
gL76UK0xAesCiFaxEJeA/Rs/ZSFLwsKxmX54LDlWDYdgCc2JUAeS+WenftxpG0aumSFpcAiqdm9m
G9F9sthl1B9H+kPMoj1TaZ+CoY6WrOHOEtF3NEmvPI4UgO+u9++UJcSDD91rgkAjA7MVkB6nNW7d
tlpMkqge48avXQCu0vNnWeLLkC/lDaCFEfrP+A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8208)
`protect data_block
wjISKAOsD78llM71QnkoEX5XUzIA8Bo4DkSRnC3tVbmfzdEIOzAElQV9NNvrdjPBxFzzGu0TJh8U
39TaMW3UxB91UD5cBVaYXxfTQPDzx98R6BKPTSnsb/CqzLq9o21j7N34LV3WcXUQXj9yhFC88TCr
YeMzL1mwj4h1HbtDKMO2+97La1bTb/R3m/KST6WzuNpY4Mh9PkGWsR8W23OPqWU0+puPySfagnCM
Zz+eiFBYTEWLJmEPGacrXwJPLTRhqYeOP1CtHPypAX3hboShEkufuA+RI862p/GrpI+ptMv9mKXK
G1wJq1yroFU8n3MiNFKxGOPgPM2Bj19hMg1SiJPGA+cnXX/v4MgWOxRWtu83/UHdbcOlBho20hev
TI745ekBXvA918jer6I8wHkXuVEHqUuXQ4rVGiUVPPukzP76WuH+T/tSLNgMmX1BiRv5e6Q6WrXa
p4PKfOjTHeAAO2ZN+dRD7ujZR0DVAvkBHFpaawQN3J5TM/FR8BRTHp32rmgCf4TjjfgutjOLjeAY
FtEOiRslXlMqVB0kfyq9H670oiUY8ZJQp79XSvw1S3UvAPslVLziyITE19tveM9yTD5ZNUlSj5SR
gdgsgWp9lNTMtfqgAyIz/WijdvJp6GXnPYeQcvYskM6ujzWP5I65F6Ou1tilSzQS2RUerxEb2MsV
JT8jCRckdkx/uIiTdMCIk3PWvXG2lsiJONRd9ZJRsDVoQsGTuJAZTj4E1HxIkVPzNO/Hg2itpYY9
F3Ne1LGBE/JhGl4t+rAMk06dk2RlAUACom9t2PTCNLNcgu3iQ1DHpEDe8l9OP1tGHGgk/sKSm0wG
cDgyw1GyogXi+eCFh6G7U4aE6a9F6bwLCN3GKjlqIbUOu/bh7ypitgYMv52IKW5d7siO4fhyiJ5u
4ZK73cXPc0zOUSQvj8HdTp7ndmUOCj/RJ38O+oyeZ+3M6WGxLwmZoJ0nOu2Kk0HLsEgNXxeaqjsn
9kIIVZ2u/+c1a1SZF4TcD+4C3aXBYBmKF6BTBl6uQpXM2ivwLNH1hGJCLdAeE3GIqGvaORpZEkQw
ZHRq68Bev7SCDOM9BjCkOf0TRWLHZEYFnKg+KTyppmG92YaiwOhxgcQHfBWQe4R8/yJcc+CZwfaM
0UtZGEAkgwbGAjBvyM0CFz4w1hDCwcgOw3HUbz5D/3dlqbwM7qk+Y/TtDk094czazKK0E3lhXYaE
dBpn3FgrULsviCpYbI4puOUrY2cm78vvmiwpKCSQs7dkcMuAVYcF0w8ccOwIKl/blqt89GFH739a
FjbxRTeKbvPD4DzJmKJTcttOaeVEpV2VCLXotH6BxU8wXojqqhJt4XXxXtfSTsAAEP6rXF4uzHBM
DGF/zhCsusJJPufqCTWhGqwYgPjzrJ1GjRLzpfIMkQxOeCzwH6823o6MhPs9nlmjoKPPKKSHIT7F
82kin/+zRh7bxoOboVbWNR0fmqRg7wPQmnEs3AtD0iW7uRBJn4lePl5QYPpTGU+g/hK42qD64Cfp
pZTEIn/9dlV+hHx9wjMMBDwPPR42kmIOYQwGYXgBkU4WKDlaHu1pbU3UC2yaU8tx9Npaas1Z1vcQ
tt2M5Guka2tSfV4cWH+b24VZ3mejxuLmrfo5wCa2IFgfBxfxzX/yA1f24AhuHqUloBGDtWhCfTkI
RSDGaOZgQ6sOpD69CyIsLnrtC7E3a4wVMqoxrVTy8EdWuKqSZYUqq/jBDegUslRxQQR+KB/go7we
8uUgWH1ZGYNOv0C9VI1IXCt+RZhDBNXEnSIIPHkCeBpD/QfqHaSg17pPlq9dAd/y/IaY8nNDs7kL
abfAkqRcUDYkkXUQ2KJ88MCGV0y4xXC0j3o5tsoTQzAFMm96xx/f1K9r7NSyJk0IyQKFz1cqrAL7
AjEj+Tu7r84rdNREMi2nuVhIxzXAG02zyvDpIv0Xbd22hb+GdnRz7auZMyFFyScBVVkZUoxlZl/J
x5fFQ7pV5k/MvgXESO45S1EG2PaBHqLHdm5v4oer7SoOmEn+4HJxxX5UZ60AySkhGzr0O6jnKjd0
2wuZW5usi+wpAeHxcXSgifRl5QfEty6DNNkU15ukxzb9nwnD+wSKzPArna1abyfmNKyGQfYqU43z
ZEpJt+me65VxrGMS9i4oR2nCXrJcJg7FbgDYb0rgJbRFb3j7zxm6iIzawX5xekE6VOcC3IK/1+xK
/PGuYsc9za4CShSTTsOZJG8yozNZlvXk8uwuYew9Wg1o1fPhVxmgWJvS9eD5FKCdokRqC4vN/45c
9HWUBt0qnR1kRgCD7sjPzHG5UvdkcLpuhenYvlsoqqMTGG99lr9Mc26UdnkTC5ka2Wj7U8udH07K
pE/SHnoZxnNM+5PpBfmVOF2KLo8lHMMgnf35jZZdcvYhHdd1ZcIVCnHfzvZh+tRkzK7Eq6BxzSzh
x+rqZQ3mLr2Pgiuh5s1yBD4D5K4TxZqxsIqAQbGQqvMEgCrHMxywei5v9bZ7tD6fy538xZclnPBJ
gLwGD4sYW/aClTyBh+99mHJSYP6NmVLwsG8j+Xsmsvl55pSATSYunOtm2laVYWiwzcR1YDJKBfUL
LhjuFU4HYV3452YBxYGTuoj+TLrSPefa1EB7TYePy/MEYgTjvkn4rTYVtlg+5ZcVFGz9+kvweCmo
8egluoEfWYDXi85ZTc0FI3tsbncm2FO5zxF+zSbhOjjFqA5navmiFT1vEk5ugu7e67/BFRlHkAfc
hWs5ZKtt+24QANcU1mXzld5xIVFIeGo5s+ZMnqe+fGi27fAUB+GPIX+IzDtsr9luBs4M2ZTABjqM
hDRROXMxngyM4q78CanFRPHdl978/kvPeTvj4XKcgYQcmVCZ/QnLnKwj5BECBNPnVVfu/tRbNBnQ
Wyji23Pc5Gz+MTMoWvIo+2pZ09Bd0tUPiH/eP3/rMweu86eD90wCaJEqR2UZ/MP62Rl8sXiCr2EJ
L00Y50tHJd3N9nnsQj7rEpfHWDZebU4qr7QWVac32pOeXaB7mB592XM86DRCCPxx4sCmsJkJr1ON
DweeLCJ7MVaUsQLZPOJH/fgaLKItDA1hkBEDOfLNSA+9QBcjvf3ZRobGq1h5wvXag1pFTrwyJdAx
zYqA3j3gnOo0+rALD1aLGRvqd5Lz6PmaU0bHK0NmaJBPsaLBco5xWW8DKflfsKjLehxGkTMclKwT
gnUFRrjv9FW3D1vbJGt7+8hvYGZa+tn+/GiT5vvr2Q+eOUEw9NkPhYhm9pAoY7bWCbf5UfAD9Cf4
sa0E1t/pZyqiQUbn9T3U5mp399a0n9y9bVgbk4kRYWPrS3l4isV+JPxSeiNVjLQjlSv9Sw+68lfY
FwQ7yhfoLyao/laqPvljRYQ0TTcSujMeIiVoAZP01IC4pHdOFCIQC0Gt5To+Xh4vna/7qzLQ/Rm1
o/nnhPWx9F75TA3eYTkmckl8UPbl3YKRGU9QZGiDXA2KdDEfZI4FXpAa2vzG4t5DugQ7ysELf8Re
Aa49Pyd2ovMYDOg21Mb0YVnPpaB/aeJMaVFv7OW2w94qppSYJE1P2VpbpgNxwlh4ak1wzpe0IvG2
vMbBdUBtND4ireWgfOfSmMMnrKhzbA2/H+KFlrhNotNk5rtssp+9uuUAykcZtxmGtbjGOSJL2Tvw
DXLuB6QudzYC51po+2A+0su2cLmRP193H9mHGBC1Z9t2CH6s+Gt/auRn88gKLzfLGJkv+rX6KKST
Qfw0whGysNXGUE99qhdiAxO7Bh6Em/4+dESEFGDdl4Rf/Y9OhMWDETneUziz5wKTwGiG2JgoNgTN
f4nNITjNhDlYdzdUfj9Bhn4aH2Lwn7aAwWzm2VwpMIS1xrhKavLPb5UQDzf2oRwTDv4k0BOravAQ
YBKPB69u9vSygAIY7xogWqE3Z62dRIYnAw9kf2snwIfbhQexBX1Js3wkLNzCmgde4+VUgAapVr/o
wpWuIU9oLpsMDfFX1vHWUib9saaC0RHnN8XrFNy913O4cxis8D13yhQzC3gVOi3AOQaZm/RPiD7d
eXpvXrPLQMtxdiKZQvfgZYlftdL7R0TwisG6wAro/W032OkYSPYShR/Cf41Zu0B2p5V8WMdbwquz
kwVRJ1LO7v6dKKP3J5suXg5LO5O6WJx+JAuDRlQJPa7hoEgsjGgUyjSoLwNsofNFl2b/sWxLVh30
wXqKfgKZjvzgQ8wtjxexHCpqxT1FWqcvag/MkLdzSDw2nFcvpUFFPEjnAQ5qzSqRpe8q5jTUKzl2
9l4NOFiXSLoBdNgGck/wVQOiQ6KiQ/5FFq5uNb4rn0Wv5HeIO4KS9c58x/t2dOKv02lVkULDoUj/
FBorlrtin4aEgFU5BMAXV3UVJOA0iPvgjXJNlzQBJLQi6KZQ6neTzC4eFUwjcmGUW6Mp1y2+suiz
6DEMa6oEkotbjmvRUJOWZl06j6lP2QeSrdf/r/wMKc3HEusTUBheVhE5MmbuxvkGhpJn9idqoavV
4p47rC0lvf6RIAya3qtFvF36XRySWZuClOxklKgnMDIjgvm0MueR7RkiOZ4S1K7guYpzZ2tMksLB
HmgOmsdVrtjncs4zOib+QonX+H4FFuxuyMwBXbDVHRIKrk1w+Y3ylO2axCKVoMI/IMjyFDnMwMLD
QOjYerWkzmnWovlCaHMqrxR6M88UtXDfZyinHpDYC42SFJJxg8d85LPwKQjUA8Qi1KxwoOK7/JR3
iWnbX3Vab399KNT65YDpppKCEWA2XNYtDhFbmzIyaI/76bWImF7nrZW8dMcVRU0oNTso+qyg9O4I
oEU1rrxQ43TAjTVwChRFHwfoTkYX2LHeGGrzaAwTRMYLs2TDxJmnnTjPP/YhRclSPo+HNivCvzI1
AzrmtBSmZByy1i01EQkuGHUKCgIWxkK+sjZUJgzpgNuyztiwkBcW5uNmKyK9IpyeMH+fPToQMPW3
fX/rlYjHG/kLUDLi4bMfwu/CfilwfomLC9987knafIF2sUSXhdRDJXv+n/CTQJ4ak0kndjNF3uvy
R7GaRoZzMIDhT1NLUNLaRAqPqmKZ/GRpNWXCNufYbnOIxmPBh9q9wmZuUoVf/ck5Hgx5pIBVL3M6
YgJaf5Bu9HW1x1k71o8RbUbR8AkGeuwwmu5/4JXKKND7VLJ9QuYpVOyigw8wBi+wRJMJbwwKTbuK
kgHV4ecZZDiir0adeZIXdYuVpIIo0SkUt7bl1U/wZ0FXc8RByWQH8Cd5yVeox4aax2AgK8g4JPCc
4deyya0lez1G0jzOsWmmUJDiWm5+1ABWRlNfGO9sIl8VIvzyvBrbPEtj5hvVz4jyWB/LmCTPzioy
gHYt0fLO5Pfc+GxY93atEyHQmjWp6Y4qBh/9BWSVPCPf6BEka45V0rGftMnJyST3J1ykuga130ZV
kYerRhwDTrnwF004CGFd7SuA31eZ09dn5uaIENPStE6Yyf4Vvlnwq+TNpgYJZdE7CoFQAa9QXoEY
KItD8bo46luL+iH/raQ50fb40fZTTl7nw3kYUTiqKkYH1V1LM3TH6U/NYHleXLsggiu89WhUFKbL
yPaIXM//oryvDRzkpCQ87Xf5nVuHoWP635WPys9nukEg6sP5AZEi3bOCkFMysADKAVO8XR6V5cdv
mXNbsVYAyXtFgb6pRqEma9MymnF1TVVQNpYrLvE1ohI8W6igJ0/fxSouuSllobOIZHWdp757mu99
zMXkt6NKQZYQTWcLiRw4KhbSOGGm6rSJMVCZS6saMKjedC3xjC8u15ZRn7GGq5FcKxOPs2bSTMdN
sgv05Rv2k7+yMzd5cqd3ITs9ESu5gZLyqUHhZQKAsMkPnu9kdHNeg1DhMC3/HmiVXaUJmFI/gxic
0Ryv7978DDsAPJyrpttphIkGoRY9D/V+kGNmtD6GG7gLftH2G8QzbNcGYmH9/DFRPkRDmPbA142B
fxZ0SycHQ2jWsI7xrcWmhb3MjlxLxyT61V73gWxS1bKtgxcZ/7a9wU/z4YqqGU4IcBXep7J1BuL5
4Nmqc0UYurNjDtvUDwCU0+bc/7HKlH8L5YIScq56ex9WwxvX66tJ234U9VFXCoOi8KieJ7cCaZMS
FzoFk5gM/eDY4pp+GJ7h6zHz0pmIjyU+v77Zzt7aNCymgvD+fXd10s8g9HIionuNhTBaDDwCmUcF
tYaXd9g1c9XPVjf1u5x3MkfDjyS/zs6YzJr+p+2ZLPUzBhN3oahKBuBAKW2fMP73S3DGsn9Z3MsJ
iBxPWodqKjFgGQqv4ztHzRfIZimRDpJzoOL8s8KzPMDnQ/WmJb6Tkrh416WJDZjZqmT+MNmocTLy
/JfTnj1+N3YFQbpEYRzFVFwUUOx0zzStzaXqHeE4GpmyGiT0oHL5qxCkrhZ6NxnNFnjBu1SURrXe
hW3WfJVmQYuMhdUGdaoNF/z1NjuP09DZK6+qny3oaV39oTwXa6DZsg0u7crw6bPRbnbgXL9P20FK
bHe0f6+Yp+facKXVZTnZBMSYAltK2NGK1y2ZjGUqt0E6m/eY/wamQqmctWS2icYhB2/+cCZlGK+K
O4WKEKrBKA+M813v35uxDp4l4SXusd1US6iHJfw6tbPR3G4RTpE1D/MToeW7W8vNj6QIGpvbUA1o
K0oFatOS7P7HCQGbJFd8MY1Y/uL7jsrbZfU72ihoFzaPqP52PzT03iLlFAljEzcbcT52/aOywUFo
tLAnLhzEgGEY8UbdWs7qlbqfHmXMuWWVd1ljM4ExByu5Ijpdi26Jk9GF0NdWSls7kBNEu667ZyzY
yXQ13d0EpBu8B65q9dYWgC0oNqIaJiDGMbD+q381LKl7XybSGJZuajFwyjskd5F31J3hoTKfYA6/
/YT+hSI/Ijo3wERi6mF68djKbPW/34ZgRN9W8UXaJHPB9OQkPTdz457D9iDiSDijHnujKzsN3nGm
s/7c5X2G9u0eJILj418uvMkva/SC2h/Gdtq+bO/niRU7VVkz7jwqIlDaXGSqP3InhDLgEArproow
g+7gxd5FSFh1a7ti/Sn4Y9oxyA/iqKzttW27S73t6QYIT/MTnXb5PeE9XxUu+j0AoXMhT13SwNRO
HS/ovz+nzo91xMC8+sntQ3VYA+y1WdAlxrUNdjhYUJuRRSVHgAYrJfAQL29uDCFzA3HWtFMO3+ee
CHT1CG6PQWBCIXJjOnjfhyd/Snvxmot+cK7MSiFcQcqLSKWpljA50hvjLnebz+S78FWb8M24Gdsx
1GgI1VlisKUyWcBgiot68M4Q1PRuiUIUjqTJLMVEhMxd7P5kvDYredmg+yJE3wf8Bt7K+ZQaoKdw
SRk/+zahs+8qfitDqukiEDDLm6/34f/h9/v+q3BHRw7JRjQfZtZ0qya8E7qEAroRgIEyZsrE3awa
ECMUgiKYKvMPE00K11EkA5xyQaOBDkKD1WNUdg/QhN5AfBE379F1HfyrK/ehGTl0xLQz/UowTpMd
FIU31YH9v3M+3/nIwrv5VVpqfwp6HWi6XlKljh2WDQwnEzzBCfoCztI312wLIlFTep26+dMuwnCN
wqmkNP7Cz/b2TOcJnxq7PXFR3YvNspAB7+A5bg3DI1o30FkJ6Jkl08+yYOqb9+axngw6oUwBBDY5
C09dA4brbtqnzBOfEhTqEUCFZnUotPzGf+wjAmyCqf/s4vdms6edqYGR1XZx7RXxn9JuCMa+iyNt
VgVuPoaEL0SnPDAd+RzaFqhFrJwJvDUttujdkMtWkENbzWvGRLM+Whhp+MLMO0Ku8MQIR0IGi9zu
BcZlE/964TP2INIM0EgqmbfA+JE7ze/sQorlR2GDo5BYj2IAfwrm6gtHYRnWD5ORhG9FMffVWyjt
lxiZiwouPUKGBB5hF8o74XcIU5PDSIEzhYYcbXtkPVJ/0bg1ccUH2Zq7AoMbE6YzV6aUTSvRXnjB
fDSjkkhJVR22nTy+nx7EAJnpT9A3vVPgLknrnb3SBDYjHChaJn6j3yw55KbGAqmzidXutwpaEMEP
RDjPG+05ut5yo7XaeSdpk3nAgvBm+Jt+y7Q2zzE7OrT9VN79XfD0MEvb2vPLEq9kT4guvF2IfEA0
EvtE4x7EfqbBsdovKsEP5eCtHve+sitUYOQvmUNqns6qtCp19LNfEaOZkN5jj0L94HHYrkWei7hw
9J5LpB1/20lR2KzlgKe8iLTQSZ2btU260pjmiKfhRrDmwcFJ3KzJw6l1DoZYO2JixfznR+C9oAKL
jgTk6icx2Ft1qXpMLoe2gcpmdGYajgWfUG4YPT5lv9hyVc0WLDIeR/E/EeEQHCUCQgsJdTQR/Po8
lHae+zh3zPv4M2pUHFRPYM2RGwF/kvyYoUWoGUwqbF7F5Qq8q2Ma+Z3oANwIzTAPqT9N7y5qoWEG
ctahDpZ53wGVq+5+TkapDJ2HNraXBw3NUOayXe/4qW85kHnRIwINfvBN3CjalZ1UwU7T6+Iyo8e8
pjlMUAjnkzrnEZNVZoPS2XW3wYUYhYQc+c1wlHE4a1mlaoEOA5GaBXTvhQJ8Xcl69C0WvJXOQmmS
VNe6pxjwqufFQuTDnciLaIihgwU6ZFwJG6K35B7japdzF1YvFlvY+Fd8XRfVByMli7jGrPiwGrOc
40lm+aPK4ZYp1CMTiAv6NeOVGBtT4E4tbaExg502Tq8a2De9JwRub/+EBYVHQO2pJ+4kx/ik/eVU
bbySUkuAPu/9KT90JgXKaFikmRR5miphJOAImqx7dGKOvHHB8jtK/wt7q1h4/7oB4swEyv08k0++
+NJMLdbcgBVZhpaqA2v2O87ghiaXBgfkjoULH95xFhFIdSXbZ2D7q6td93MTt5XU0YHn3lDLWfjj
Lc9HUnqMmBEgOrfmPxVyIqttE893HW3CphQlildYlZLP08vozkyP51RS1YQAHY+qdEgXypCsJSgh
yGzISW4GNYe76ougXAYMJL0Xb4c60loGsP92tkLRMzis5VE+Z0L+x98ytMY0cTaap69t/BcW8wwt
uvPba1TaXLSk0JMIlzTvQU3cAbO58wCMFHtCIEVyXQ3p2kxTxdSVTajLlRHPzttfWBpJJdNXQRAT
9r0mShyCSll7HcFFl/ad+OxsCOt/qvon0O8g2ti+EisXsgiTIBiSq52UnafPHRJSMfG/STzjtLft
T/UJd1I/6lx/9dp0rkGQk4aar3VIyF80xLFPyxrLRh/wvQH11xy4YuKlof4bb8jSMjjPPSOrulbW
/4+X8DKAPYis1nWmWdsaM0mAs+1ubPhDt5dukCseZfSy89Vqy1+Gl52DHk3PSQa0bmQIa1Dn2id+
pf4I459BrLXDCWYvstMpNbCjnGWvu60IZ9IDEULW2oW4jGtQee1L3kWuCqsscvsCai9zELZLoVRD
OMmQDgNWBwCHx1krnnorTlvPXU4DXz9Yt5WqXkzc40KSlQdcrgF9K8Q+myaQowVS5uodoRBJiuTq
3KIogIRGDPV5ZxEwflkszq963xfF64wzKXcAlr5vfyOXg7RnVkKd7Pw/6bTWG+Fbx9L3HeKg1yrY
nOZM+65wDJ+HXYh0rFT+9EB2MZTUkV5WxWLTpnpfmG9onhSuQ8ERuwm6j06F38Lxv0QR4TqApF1m
r80AwYx2sFNr1QxC44L0xkNpqut9YcNzT1C0OGjY0w/ATKyf5Sp5lAM5fdqt9R2xW/OgjgHCCqGU
nWAaa9ylf0WE+X3k6xfo1ENVL6wkoHBw50sTIC6lW+FyMq0Us5UkbLcFmmZyvSi3rSiVnCJej5vw
jkcHa+t3VTQtry6VqSTEqzKrcSJvhtdZeAmfTjHqsJuW3KZfZkcyuilejIZCYGv5sFcgRiGuOAer
fdQNMdviO+1fRUa/uIsKJma0ke5JOAKS1qxUbgiGwTvc9CGOJgj/ep4gewjapZQqu9M3X328MOgz
Zijd6jOgmDnX30kRFbsoH63whMVp+bHt95DSxILNiDe1rlc47wp0mP0tSEkuS24qV+hYSjE2G/iF
BQj4N2IqmHqjOmMMhtxUhhaJxXUA07jT04qt7AdSbejh7I9F8piNocX6uQz70vLZYTc0SF5jju/x
mC9ZHs6zVUydw0oDIg3pu3U75s82nKixGbPECfq3Hu74N0AqWjd3KRTKEpKI3TSXpwXUfzkccKU4
HLBW3tb0yZMmI+oKJ0+Xx2kR110OxRLPcb2reBrJCGNDQGl8wCE960X4M2Uj47PtVqzKXTXZ3SG1
ywOxvtPWaCuOfOFvMjpdrlpW0lYeXKH4vQH3wU1Audl8pR89ddvi+4MtXi8ZKYxPPcUL0r0JHiG4
6mXikH51xGHgyAT6ISfs7wUHJ1MtklRDIRN8KYqKDbWRYYfjdH1AzCimPwc6IxHcApihD6Y6gNF+
+ewrXM6RRg6Io01YqhU8prNLCHWs6uC4c3IxjIaHrxlvSqI1BmaKr1WSt2QQk1Ov+ogrDW/u2j0v
MXsEK+7qTL9guQTmRSQUFEeaIVUlixozXFRqAKD25Vp8dyijX932eZFQE7eEdPYQmZ8j8iAFPpwm
x7I2GQvjH15xQyoMqTNRex9CzMfI+g+X/LOIpnL0mVu1PiA0vYzFFuS6F5qPGdFDt8dOBdDgkVH2
ElbrgJOnWHyjQ/uqhKv537u6iDQH6ZXRVMByNrkfVtgUTWa1Jt7Qge6KaIITBjYgTe613D9wrJNc
3zRxaFFxA7zgh53+Zh61iTb/M2MtSc6j9jZCy8JglOYSLdSaq0XlA39mvjIDYLm4tWeoxk6iwzjd
owz4gNDxYzXEjlsJUlj53KE1CVyPrY3aMyoecy7zhcjEOzICsRKFjvbYkPMhHtNzAGQITi0Ca8la
7mUPXR6DzBJH6LaLYPslppT8XY7xEAvJ6CZKzBxnkjrhDUmYcRppSmcI9tLgdm04DWePnH7UfqK2
IIQ9t1dgiox95A+8j+R3MTBKxTDTxp5P17gISK5Hw/Bkg/kV8+AP+OcRgs0/fvjyL+grb53GrS+S
`protect end_protected
