-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
PMcio3cWNaMCWLGwDSLMCnjffy6cMygFYrc5c/L7CUvTJ2MiUkIxJ9svxBMhSUUPqm9NoyVtFmT8
zOLJ8w6MkglkHHnWu+zqHNSyY4Tn8l0OsdZW4qfn5A5d8nMihHDj2/i2JVZ0tz29h3hOr+51ZURP
SCoUBeDH89dzxLOIS8TXFxUizBz6yWJU7iuK+/nvALG7d5305ETN89rdo1tBxQs/mpfz0Bqj8cxs
r+3lfhaRLfZ2EYfxs+KwrzIFpzHT4GA8vxRgnFag4q7IG3C9esG+KMMR3fYznH01CQwdPn3cpc8q
o2swyj13+32yf/4xOhd/JDoOmZziAKxMJopKWQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 23248)
`protect data_block
nG+Hd9LhUt4iXZ0ZX1NGofIRjXd73WybZmf/DljxQ9EA6S4v/eJjge07Yalb+EBBqq8ZoORZFTPm
fI0fjxUcsEQV/P79onow2eD2PMPtjNwyx/38mSK8pu1WtprjYKL+dzNWwVT8PSm8wM5az53ttjvC
/foCdJAhU3oOBWaxZL/S3EVBU77DA5eR0YXYkKj6D8YPOjb/TW+KvYp8ykQIltH6ZMUkt16UUCgB
335TTVjma7UGl3pvhvRDffjUNLthDgYp7Mrd+kq5pjdjcyLWAI/auIYNqRBJQobWUa5QRJHlCEN8
kHalM5n7It//6osrZQ9B8r5kIYD0FpLlqFz6RsAsp9EQUcDqLyFH2CkfyeyYBRIvLRNdtb1HqAzS
9G00HzcG9G7xAiJO9vF1IOPphdwe6Kgn1dKPYHKNX+jTKJkf+oNOttUcYdfoTDT9VQZW2S+e+Aro
v0Nj6OmgT9Ch01iO/r/2ZuLUqFXSpQGz6OAELsbUhqzGYClLnyGRao7j7gPJk24+plyk7qMOgzE2
neNblh5MinOnpMkPX1IZ3DxsPJuWjrW3Ky2x+hVKd7fedkhGW98RrC0x2WnSp50rVUxZvggxoh6g
3OOHa/oc4AXNPJwp+jKd4l2oHAk3Rn+f3NhMUVylnCvpiyj+zqmW0yvBHeKbEnjp5z86Ue3dn4Je
cyOhebvYCoAQnnG1uc/VprjuvHuYcfU0i1ujEQPGZv+w5F2e6V9NsF8VTxC8mq+H5XmipQY2ulY8
aW4uk+cgltuaw2DSNOGJy/iqFm6Ceai/Cw9oJFmYu6rTQteH38OjFerpZEO/a67ELzgeZLyrNj+H
jR/+aQZ/JAL9Ub393oVsYUqAiuOmaO3zbcxOTrqpL8X3nPh2DRTnf19TUVAnPELnDS08Gdu6MI/N
5doSqIVYpUKDegvCpyLbcD0YQ8cMBrfzvDjbtJYVy59LLpi6kKuIiSDFd532xgPrnzruVbE5CkNi
dPenIOMF0kDV8MOLfmEvqqOl2BvMub39vd2t13By1CBUmCfXSOylq9BgXuFTWH20MT5sK8tS8gOw
nLl0xJj31CYueAGWRVtdHGqH/Is9YclC3fGAv/PaG/jyLHfwRK937GFJAbA+L5D50Jq/pWghBzkF
L7UwMUZfrSBhKDpp82aIl2lWe81rL09oLQuDXJlVWHJrmAFOu2zquBVa4MnvbO3NmZZAnfV88fBO
lGAyhtgTMVR/709zm5yAwphbxLyUw24QD5pj6yLPtRDuiLBMcyDKztWoAYjc1xgTr3SVSPbsFvIl
BKHg5mAOf4gMSx18LBUnI+j0EnM3l8iJUFs1S33yc8kDwXX98xrKDPLtCCcCCKOGiLuW6DJzk+hF
+EWY7cTkHDmaapIlRTScVoWh8g2oqxQbcgfplEoqV+5s7iNJhnybXErkCEzLZQ+fwsgmLCzU8bQz
iosESIQ/X+vaIfnAS0CgMbY2oYVCFZOVWiWR2a4aJywUxvUWhI9Jgy8hYT0E9YpH1S/ucXdjpM1s
OijEbB5jGjbLZpN3WfTzAJzRdCT6f3tWwvXG1wS4R2tDJhgRJ4JeX0xwrX/MjKVR3TFq+JAKb1lT
FtJZrioIgjdm4W3mrECtHl9Y2zp3laLW7cDXNYRBVugjrInPhdjWsRp+6XGtZZN3/ccTbHCnH0HZ
3G/6KdB4ZMuOXz5w+6qzsi729qhw0i0lUYf6SG4SVQ6wsjc6WDg0DC2IAiid13Nun6NcNjIPBjrX
H/lkykq7LtHwK5W2SkWxZoj0qUeO9wzwcH5AZ96MQK9T+yBITsaBuu7qt5/Ts/M9/ApfbApxZzg/
KbaybvlO2Jo3AdVKRgLriqfiSr9Kmh1//lZhncAzESpx5pbX225GzM7S5r39qPNbPbCJzHl32KJb
VwEgoSMnvjGDjaeIlkAKuh2K7KVjemNskCjOHW5w3nicUOakbtr2XbwNc/coB2S+BylEYM6DJOZ3
UVvKKZY1vooIURNJ4LFVmRzPI8S/Qv0BxheyvMXAc4qaCY1WJvtTICsFKKf3nd47xFdhgrv3poD5
MeXPDFMIScqR/HYNdjKQPCi7/EM0hWod1BECyvTljT7G0fwoUgkm0hZcFAe0y1rExaE7JFDxu/AN
HXBwr3T7o9qnSnfS0Wo9/oFEuzAX/bCAdKh6PuBNWof7TgcFJbCTwWeVa/ndjfQqtBZeI6FJb1Ke
9TC5O53S8My61XdY0UzFIkAJTuX/MN1+iObZ7gOw3j33+p5PgncR8C1aC1/NplppkHXnNJ+UKn6M
32j8D1zPtHl21Jw8pLJBC3reWLKfPhFw/csb3g2+GiixW3h+ugjxW2+z/WD3WoFl5imiId8kwBxS
BBa6G5rY9kIGmULqKtIihs2IXsHSrI5KXvE5qWiIh1nwLkfbIgFjZaaoVtx+Ag1u3/VzrT8afYvc
SATDJIj6qmOH9W2XqFWhP7Il3o0uDZ9MhestSiUws31C5A3ytm/yTF2xLrYRwYHd0AKiM6lxEA5e
rCtSvzWMcDwLAGunqQmr10EKSbVGK5DbnS5pBVomDiHO6P6RuwZhrmD2LO0DLOQ4mYPzjmHr2O7g
CZIKEXf1FxgZxPOFzdHOL5nJqhOLfHwjuxUw3HFYrVe0oSL4vnW6D1vP4yxK4XecWzWK27gh2z3D
PPAtOXWJfC6eJ5+GSz7rWCinj2aGolcx/1xnvD/axN3tf7Hk9VzPq3wEJ+uR93133udjHwtg+qq6
l5ByfUCEgkCJ/UmaEH0R4hYz2pHkDO96FxO8j2ir7EcIF5NJOVxzAHp5ijdvb5i3HBeA8k85CqcV
oo4PP9owsGvzeUdeeJXTzqkUodOPODsOnnxLZEJJOvgZSx/QTmF6bcbgOgygZnV4F+zL9C71wQVg
veWkgRC0p5IdutxU5G0XfuAb/aoP6oSJ7P0HQbWGQEXpUZT0BTfMrvIzvuHagHcIUhnjjVuI24DM
WWEns5GSgLDy7q4w5HKrxPYEJSzcC7FyASUeMMN5sNbbAE67eaDTwvTvrDwfvmtporp8nW/ML/PA
krwsQ1qBpKKneCIWffwbgWimLKK6Ho3QXf7/TElcgZzuIgQX1Sw/qlHa//Nh6fQOy12ZFIvOznlF
Mw4Z+DxT7c3niUuoB3ZDfwypVtWDYefP1N2aeLlest9z9hQSXFQzAHQ4L5PWaOgzaTXqMFx5Q0DI
T2sXoA4cTRbl8cS+kdAItZ9hPn1miS1CGTWnEnm74v2OOSY9gKXUc2nkc40GVZ+OyXBQzXrj0xws
gerLnqIZa8QELaGDZWZ5fs4gUFgYFqgGMsBfarWtuq1evUeh77q1XPIuoRhQUfy1R07Zrnv95vzM
HwBvTqmfRRkw5bHWIKptAsaoK8tCy2AbwfMG7ifqr4KS1D6UQAU4TrEzRBHHvPtczWxcnZoe1Igw
DyGxjLX+bag+IWpcnK4uZj/NFjFMjIAILyoxnBnlJRZovLyzw7MOv3up68mip1/s6rBNCzEImU/t
jCRXZBOlznpg0EpUJYjGjj1fN0CL2AoIBRbm2hXl1Ixvzz0BV77Ldx2qoK1dtWstDDiQUsiB0kwS
oJmJYFIVuLR9m8A3NDMfGfystHJGwDnkYOUVGFVRgtlN2khD+1F4mN1h9NS7/lJNQM7H01Cat8gy
Nwg+CvbkwEg+kymXwZL1zb/KMCjapTGW94RMF7HkoGoIQO7y4xn9FreSlNbWZmUoyesXGDOUIUYe
pYVafL+UXAjyCIhytBwXHXdJJV8/R6DqggmB60Nu5ODKTPKMoEGMN8j5kvoWzjQagwSEFjduwxup
+3zOSfkBWGMR3oMvlsWoSDaSyYXFdAcOybCyq1zgp/F0UsbLyPnqQVut78mx3wJiFk2hLCrn/GOG
hQ9f4xLevGd3f+U0UX2cVnaoZmoWMnQ0Gig3d3jexwrmnki6Zo5p559qs4NREj3/mHF2Pqc4fgsW
CFnF68FPp7GTmwqCN9R4cqZ81D4hAUvtsBuQh2XFLe9mQn+Nq4oYCGB/2zOIJzi3OBKUJoQT6RFt
O9Yim/VvVr4vvnoF5AipWleqRpogcjr/ZwcXPuU0CF/O9eyb7QDBp6jqjkZiPYw3ykWCE1Jz28/Q
ApvEjbbzkaz+ctT7t12uVwTNEJpHA4XUNM/ZEpYLc054+gvYGn+gRVmECPcfOOMKiUcZMdFFUU7I
kf2ia2rHTm6lZR4U40FzDAVtGfhKxG7Dkl2QhZs2fUmG63fl8MYQwBLm7bYrXg/g6SijfkkB6vL+
hgOzjAochjSPWLulBsMcQUp5M/LX4/n/4FT65IlLSWCFzRW7v3SdwKOrYd22IkLAUNwrGSlgdL1b
U91I7dli4swUi5vh3lRPjwo19a9wdmbweawBjr+plry8DmTLpMCT+ekbRgUd6tPph4IE9jSw18qh
8Jtkednl3yMmOvboFLfa22WREEP9po9FnrufYAyof9XJkBpQchaDhzlfA1FMedQmPbrSRaIqmhDO
3jPkj5g7C4t/tHXJWba+e18HgPf1Navl3Wr2RzJFn2anI8qWJp4f1VaW2C2DnW6rVoj7eI0y72rv
IEEkFzmyCG7ilulVmWwyjF1aVzlx+mQF964qc+Mdkt3tJlzoIhdCGmrcqjpZ6S67EIgFuTLrkmTc
Jh5kkxQ7sBYXxRiD6y6pJdnOxOzATFTnZA86pjay1yKxhBKKKMxWKekiEZBmQyg2Q7HgWD54kw9G
mb9UVeNWueNJ1lm7Zwrtjss2D/Gf9rfB8Z08flH/9Ubz86kiPWSVqyMlqwwhnN5ZD62uN6OET7Vv
0LOBmbp3ekMIIJrqNHdQvPYjCs/CCvoAwX6cZa263VkJ/6Zv8ADQffJCw0zqbU6a4O5tShxJvMps
/+m804QcB6uTXMW9CNcvbgMbhLFvZtfJs4Rl+9ujo+4TNC30w1Wog+FT6vTBXS7Xtw5DtQ93frsR
9jpOwPUS97cCCFtFNw1bquy5fsClG3j45Be9wKkZY0wHtIwF5PSUhA9TOc1TTkSwP9RFs8KzRVWY
nZegSc5IjoCr+CsOgG9awQWKYzugXD1iJqhp05Hmxc82s6I/TpKnXasHTCM3Q/Ib22WaBSmVJLhA
CV87WEd+op12HgEgIqN7pYiEHVQK/txm8VDnThBcUnwLo2SCMpI+S8qGFP0TAVw85mUl3MQckvIK
kylc2QzNs84tg8Jkbg8Fxm/V1ywqwp0ATVTeVs/NFrjl4sJ4Q/63wOfOre8IRRBR/r+LzeKwY3+Z
OoDvKHcxVyEsIYSNjG+UulpSfCughpzbmsb1uhnc4zHK8jLddLZBp4YOCr0/nwW8ORnLX8zvky37
HGmmyZiCk9MinuyQ2p6eUDQz9Jg3eRizWUgQNAhodMU+Y4/PEh4fWuK1jSKHs/ULPo2VYxvYQgc+
zeExVdPvoVLvJm2Grrae2y/8UTZeaFLaBrHjtb55tYwkQXJ/32e2WWV2dtkzuCZgAV1Pmh+qLAIg
8WJpwfiUXT86pxyPRBUgCC83Fq/vOxb4czutQvzrBIJfrOKXdh1HA7G0LO9c6ODzzRd8+QfvLa/q
+3WQ2ltABrKdOXAX7SmC1EO4EyBRl1ojOPV08bQBWpnepsd8lwT/VeuUidTo4yxoOpILH00tuX6P
RGlaRnxvcGH7MI4HAbSH4gyR2Y8AUKotamJkQL96wOzjJkxfWzqdhJ8Niwyqv1np2XO7RmuGiQqV
NKRO5CFIYwtcdGDs4I2Jyd2ZhD+h9YdzbEYoG9bWYR23D/Q/3/gw3cCQHLyWvMAffPvCpiGybZn2
Swoj8PWBz3m6AUQA4WsWyScwV+YK1sKOf6xcUsOJ1039vZ1B73h4OAy2kfj2pwumQgkLp6ibSMkc
yuh45T550Md6wl5Ig03pRH40JbmGqL7vGZHDvvQ91kXRgBVXdC60ELGc9fwFVjmCIVCNN3gSdqrp
d/gWUa6O1KMX2orm1qd4Nl6cbChxXYY9MwyHbSAubKbBmnMoj4Q7FFWpMJXVfmL2pqbYfT1/c6LR
Unf3W5/BwEj0IY8Pq6Bqo2PPRbfx+ULNLJ8NY3wuS0u1kymG2hZQ7c7ty62IMMH66XrmbuaspvLv
pthEPQfxbtM7/tmw5xtSZrDRtYX0yyt4/mUwWTTjTPyjWmYvuTiHiLKnfwRjFNKvkm+oTyWkVmO1
LAlXDVnHJIgaAz1uquRk9hoHF2iTsYuBOXtZqXaffKvfDQo8Eqo94y2Z/uIu3hVdDdW3d8w0YNsk
/std/4pQt4VwUNBVWRG9aWjSRsjI6ESidfwMTSGejj4NvArZudCqRJar4eFFpMnJ/A9hpBvLxHuJ
KBoY/833FWhPX9UnbFiAQ9RkYBnZaQSYYKZDouAN5IrPunO3uSNR+0xKKeTvmoJsDj5RK0sVhBir
UD4IpNcjTienwhAZlI7tCRmcaOvKu0pinRha3nHCPzzcFJkcppJReZaDo5QEAYkOfdu/b75LQl9C
PnY51GDB54McOcbAtvdFPIF9w6a/5TFyTSq1CJnxhYPZDFW1wGuP+2l+RivyjZ8XB8YEJI+wVeI6
Xzje1l7c/qboFOxGy9Kx5MrnjTY3Tx8H4uE5ElOWBmG3p1qt09coBnYLXfGf6fwzvOBOdYC2F7yy
t709sDwfTN3z2lNuAuyBoNaz6JYTwNHE275fwcbUkazjoug+bra7AhIaKlUNfv/bV7xoRM8Lbp9L
DIiS/1uBzkyeRHAwkekFB031ZQZsJNsACSFRXPmAAwveTZ84a8qunSf9H+Riroi0E0OgTe2xp5D2
2f0CjPheVESay7FrwW7Pnx00wcvnVUSdgI7SKsmEMpTCQM72f6hEMyja1nSi+H3UisQbn2kva0/G
CDQKHoU/fAO3z6aXt5gJw4dbg0+gfpolIFCd02UNb6sjWSRBq0/p/IjsFM943V9aDO63bw8mDcn5
cpf6F6bVNelwZvB0O5EEEHWd4HiLdVRkNoPI+5B11ggt5nsc+MYNe1Hx06xnmxnTOY43Zi8eSYlu
WvEK8deIyVRqxkmecvwwyLcvWRoxuq2R7l4EwZh4bwXp56Ttrq9TM/PVosG3pKyzHcwdFU3S8yMo
8I0i5DNRUGrZ4VwnBo/u0OwyI0RIJmuqCMSG/4OVNKMZc63YlWQFVtNJGGbco3g+bKK0kTcyw/iM
16Qn7HEHmqjYiAWqjHPva0Q9sXUZkcYVJlAlW3MN8i2WJfP/0IerDiRvA/Ja+KeaNcWk0AaUj44q
FmpkNr2B6bLgtId9ITLPVrevUeOgvpJRulaoVrLYHfZPGBYt4p2A6swku8ZaU7R3LeOTqZTmWdYA
Kequ6mN7SdkW7thx0ApaVj39UWNUsEjXZRN0eRe9sbp01HTRf67rVk4cnKJp/Uy3lRbHG3Hs+Vew
LYGrQpswlA/FLJEoZ+Etx4JlxxBrBNszrVuZCgA3nmJcVjZDLQW7huUFYBwxdTB1azq2TzWoV7aa
BAflCdQSYLRFD4hvEMX8eF8rVkv32tBpxSCe6Kysei0QR6VK8oMGiaq4yhBoozebwtlntQvt8fDi
MeXYmX1greCT6TZZhzMyolEtZPQYVMr7dIbM/3HVNt8zf6vc8rFxi/Tf8+VuBNE5r+ipcdZcyKBC
5fmtLZdz2kDSQ/Yzai9YNXOMeaA3DwG0kawdNh/qp6JEn8GgjYHvZ03UrBJhD6e6i2hyYX9PaIto
bgi2Tla1YUaNh22rr8ie5iTxO8zPZ74J8I1KDKHbn3wcM3lQjlsspDcG0NvGRZDtKwXSuSTpMJ3i
mrAwpG4QuAUbGTiETRgV9D6vIwZ3QFDVlxwTsw1pNPY2w044K/ObfJzbBnQejYoHjcMq988eYRp0
dNWP/fTab9klkPIO6V2pqLb/PJeZyr3Tbwqpq8MlltsENrMtbFVC4iDcC8b7khjuPKYUaWj9lYdH
LyoLZQ0MfgaGa0KQOuiIMwAQFvzrpKFS8UTi7dnYdYa46ljbT37U4tXxCJ6VnFoWKLxckjjEy8Bu
UgG0Ofea7z0nFw4xJe+1rOjxyL5Xu8vQi/BsbUuscUE4noPKc5Jy4dD087H6v3+5P2+qnxIDMnEU
AQ7bBGJuc/Es/zgRPTi6QsifFazdqK5rx4/vAF/NjqZW3/AezYAwfrpgUrpUJxv0HP5Q9Jlz6/gf
wKs0vzsHQwJloJYrB0S0gAeZEWcDTH92cittD3g7dWv/qaCBntyyTelUkBWujr6I6v/q6E6khL4/
NefIE+H1zRN+lNh3jpmR36V8RoEJUf72uhjLLq1OfcmrepVzr2uhvQy26uMli1iEqtCWnwJNxESM
rblG1zNrXafvOG2LCrrnwZJicLfyPk4Qf5aOfJ/igTtsU7Ppxzr2z2HttpGXSAhNERLVOIH7lS08
bjgZI/Swjp72cqqVRtBgGXE8ItJJ1rBst1JU9H0vNr85vKfdUMzSh/1kBw7I+pbVtuGHWYS5JNUX
4CpQR+aXVbo7/dYSCFp+92JzbtnuRa2K2eOVBr8ajXcJDrBI1LARtHqVhvWlsg0FIP9RU+LHopIz
pkCIG+Lw/AoHTF7xPPmssS3EKFdG6xqRqZBlWdf+agxowPE13BRlc5T6th+T79cHAhYzZMJZ0o27
RXjffjDJKYvDfUwSlaqoBqdgEW+OFv59tqBbKxjyYWO+6BzKN7Fs5kmDR14ZtT3ySnxNVMRZH3kK
d9c4DXVldfxZRSetAC6JSGE5YW9FjJW0rWJ9XI2vlgN3wrH6KTUdRd3wGVASuMZBHmeWQUT/TJGr
HrAFOagACEneEmfNt2loBBPNQBpLUiSFOUcTJxRPpnSGv7+mLQGx8YxfxhjkwGMB7ix/TWWUaqUC
3qm9jH0Cd8uA0BDOoRCz9zq3W1OgsMzmSjyxCQLfnRq4fvfxgPQj2J78ISqJZS1TbTuJg7Nw9f/x
rPNsothBVQoRPZCJCxkarm69A5UDmNTxtE+2RnYxqSCHfDo8yfLOcxOxvXD7EerZG51JaBkXS+k/
xBkWI8JEBl8nqdir81vdcuEa+3ktQ/ZK70rcT74+8vfUYx5De/JsTta82/vSUqxRGhpEJ91agtz0
COJhbx6JSLYmN+UXmz1Uyf6ynQmHLwYJ1Q4/AoQxHkIo9PSkJRXgrp3Yz7ZGtOWSQ01nWJvoopdd
6+In8ar0EVFKPmJpoWcXbyDmEvkLJK0I9UW76E10A+xouuaEW9hb9+2jtLLsJD9hGQBxLEw1Hxno
cSFwDv7mxQ9xg3fewZMCSQe7lYOqboxWY9eXd19qirJqpN4kfxwKuKktE+X14vR1LGj+tGAcH7y0
vkO9LOOkVamI6UYROgDPLo2B+e9tJw0W+YSqeOuVeRYP4euWokLmGjNsAiuF7eCILHGCat9yi15h
bdwV4VCUJD0WlqYhyukL7UFJ7z4JSS065kdZ3ZqNfaKpvDlUakMvjlxPX3tgdjh/AugAUo/g3Rb+
HjjglljZTZch6Sa6CGsti4nsLV1vB+tPWhoyOg6itfzEPdvfCzDayJ0k3jTl/ItcAsF4E8o8yW2W
qODufktEpFqu2vSuucp5ZaeGJHwJru7xcDqJWRWnX6D1rfwBIgv/O/Jcw4MX4Nx7yyZM5LatIres
XeiOS9e1WR+xLzhV85mczdfU2DEhuUSA9x6irFu4oEK2appG9pFO47ESwSJMhFTNVUgbsSOfQkCA
HX1/NhjaZ5a/TjqG8iRN5dvDac1O7sj11LgmSeNJgWiGrGob27DBwQzZoQaZupZUWp2z1WYZBXxR
QB/5+ICx1NujkbzEWgbFC5lZNNU2JLcaYVnmzoqZtCeWEc45xcETMdq7BuWBr3HyDtgZuDQIJFhE
Z83eXdWwg68Nua6DXxKRtjjMSwWrU4vAPONA5lSQeP2gWGF2llZS5Uu+P5PyL0mGrxxLV38AiKNk
UOAqnV+oPd1uec7frpIjWmBF6C8M7kOwhAGx4z+y4bymcXs068ZpbI/Q0BpZ4qSzQiTnKqVxuKvc
+MsLb40IN34chcH7yu6mVP86pnYqVAp32koLg9kWOjnJ5KgyrWJEaf9uxnq9B5doUAALJUDIHoAQ
spx0DHdvboNNN0B5FOcO/tPuhNOvnhXWl8nQhgsg5DmmZWuLFtIz8+qMGKvNOzkq51CNElyN40O1
RUShAb6xag0BJdOHatUX8OvOQ5d0kW3C+GWKztTMWggkV8uMDkMx6FKm4WQa0mlnA5Ib4kiUPF/t
aR9yJu0lvCUxxfutC1HiAFaXjdZLsh5yE9oy/mhE3r/EdqXF/YjV0PBluIhfRUkJCBRTBYfDNQdn
ra/vWdfOrqm6urmmxjyi+N9zgdUazflnKZ3Ugdwc9Qfc6gIRDUFKuaQwDh3Pycsxembsy5xHjM6g
iu1Pv1qmMhk/7VCiHW/zoZQZIN4GHpFKxzKSn8cnuanP3RMh4H64j0JINcPzvKx8/34zYdcD2IRb
8oh7GdOUbbfgmnVnRQaFUxYkjKzjB0x0T6EklAZ37UZXRBXbhEIySbwV7bfMVFWfhVSHgSc0cAMq
n9cVWaOCzNq1qGaies8vMq7CzJ9uhmiHWc+QFjH4H5S8U3A0ixB0BREdsuj4WVkIY8fz3INWpPbn
F37QgACy32GNda+rqJcrRDNq7AqyLxa76fO0Ni4uk8Mx/R6SqlsTtHXpgcL0ZYg+/ukqm0QTqXP4
yULrJkeQXZ68lwYkHVl9WidILEP8fJCme/FfR61q9EigBuYiUL0F9YTFQkYQ0L7jxeqtMlyMq/ZG
2DinIl4Cn4FzRXrXYskwkvJjoJC5f0Fbjisz9MNNJVlel/Rj9MwXr6HvjB2vPxW2c5+MzE5wdF+4
t7RtZ1GK+wpKBMXQHMvVeCXS4Wa1M+xKTm/w0R0gAtGTkFGls+X4vF2nwMlUgPYjDF0sNBXz1twp
bmZqgWrBTsuinWT0SB0GOCZay8VJgLvO/kkeKspPTIK4EmHnrNa2gBAQig3aI3qySNM/g8AyxqaB
4orv0IF3Ar/6D/y7l8TbfdZ+cvCdyjFmgCewAAGQLhAPSjelC8Qb/zIKB2TtyHTVHEW33dihsnN6
9zIVssFLIvcD3AcohtbPRSBi3L6ov93TbggOQRWeuFR8RC4uAeKiqleA22kzf3Z0bK53p3FsN7+0
DO0Xk9Zn54pzFO9FEBgW7Cn+0zSUwznPeOd+kLKdQNpzcVjCXVydvuOo9FxSQQp1lEfcEcJOo7I/
vMgmttxSMNKueZCcpY5Iu7sQruaw1OAx18FgiaoWaSstMgqjk0JbJMWNkGPhll0GFyfpbvXTAN7q
BD0fpVyHDXLuO8ZZgo6HiX9ZSVgi/TU9tCU5oKqV4TJpSWqPNnfkovkKKaxIzIjX7CwKBjRqzs34
RtzVwZVNxGCMX6AGNu5oBUPuZFJaPixfDCOGX9Qx6QFTTxw8A3QywXHEcty6tXTJ0bQWFWDJSF8n
cIhPlove9FwY/k1hjckCkuqOZEkTwlbUpBe4dihSDjnuaT+jbHCuiAPLDtlQuq+J6ZiuoRWDM+SM
E6iBX8lPoKLsnOLssuTQV89QjaOnWbQJkX/dcpFq05e8ZqeVFqNJM/2e8jx+Qp1gSSiaetkb/rBD
rkmotRBrze0uFwXZyJ9EmHRL/MKIaBl6g69M2pcVw4h8mlDMll1qQQKdKPi4QkcKYiokgrV7JNQc
RSyZk6Koxoego28XCRPx+1lSqlAA4T8Mqvyv7TrkcBczGuiEJM/Bad6/nwy4ID1HcKQHkJf3M8FH
v1fCaNpA4GSueEwC4n1znm32itR0A7ZbcrpHaB8hpRr50OJdZXoHxgU4GK92h2eSoFmzGgeuU48y
m/gWEb0DEijF4Z92O9MWVh4vjyPipCshPmujZq0mV6oDlWJseBiFbw0/5P3UP7L4hDHH3eqyHJ0I
rGgiBdHZbNtgOdVEG/I0MJVf6i+5pKwNkrn+R7a1Mfz5j2LGhqsHLdruF+yjrHPbG9zbsPJ0MDqn
bVY9LmiPFqf6CKwPkmj1COD0jIjq2izax9n1ixJUiTijsaIE8bY0w1VxLSd2KCjAuVsOx41va7O7
7OH+Z9mTRI+9bSQn+6/F5pTtf25Tk+IMehu5bZa7A8q8Zp27o2Upy6PljnA1bCj2RbMSjtq8vFbB
kzgBOJIrIjRKcIx4K9FEtNFzRI60NnOec/pKGhfV3naRg0XhIH/0Zk+9pwx+dFBX1lIxqOI3VFJu
60XSq1Nu3IOpTPV0O83OlqUvhz9PJxq1MwxjkmymcJwnbJNU31VoqXH0BeYFDRoJ1lryuGFsZ0SC
gVupIo2MnHhiGDvFn89M3FVsjXarfj3ybsaXSoVt/sV9EVK+vvJxKzDB7s0SeC75/O/FtcwWvU9V
VvdV5A8hTYo0nF/WrSmwwPEXHm/vDdSz6U77Iln393vF9JoR9fr4BNfYW9kJ7ObYLKjPi13Hz2u1
KqApPxOLVeE5bQYEVf3awchZOAdH9BfnkNH7m0fe+0I1G33C4GS76GLPpHAN1BPp68UzCU9G+C88
+W0pcUrc+vxCcm6T3ucI24dJzYA5REfKeJUNgEYILic6YYfvQT2fo3u4R4P0fZd8VWiNcO+ciY1i
TYpjZOKRybgGCXbB4w9eFm4ExH4wbuAdI54lge91yl/Mo6+p5OEBoiy0R6m18ejlZDS66QkYfFS0
x2feaZy8UCudvxHNwZlsc8R5jHexsOi9zKAJlpmnt+FtUo5nJ4LSQGnrr/rRf1S9j5zFmf+QiRYp
JrI8YkeNUm6504UUgxEg66UdrUGdih3xKpwFgdVnjiojg78zHrcTt2sJ4VlSrUvVNCA5kOa73Xca
0Xy/fdYitFcqjlfcSm9B2wGRIJbofLdiO4Eim6WCEgyxA+3Skp6AaEgCfKJxgib+bZR3wpApYxdD
9YrzuHBnr33SQOAWiP7hjP/AoUxiHhLKmQ3uLeTjwhmQ4IDZnfsryc0WWBuaygtCl0jluYggPx5D
N6ZPbsrU0qLOkqBhi040eBEevCNXuv49R6H+9l1+kTadtfYwq2vZp7GFDOEiz3lWUMdS0zoADOh7
wS+HaA2fRyLxAjEfJVJrWxolVo82bZwdyA9c8rpu6vVqW4FOaMV88DQkZf3qT5CWXSS78uFzpRVv
2gpz4RFLkll/HIO5oxlc24g7NRmmklxp4U1HF/uCz6x25Qz2gOTkNWUU7fB9uSdSOhJ07M6PvAQZ
+Uy4fSv/+kdBBwIRHQPaAA0lAkO5G39oJkBocjq7/u8XdaKRZr5Sj2Z3Gu5iGdUEM5xSrva7E5h+
4DbQ/bz2umTQ1SsOg0XPLF/eWIcQVYwNvvQCdSvRNGuckQfTBhIqzUv2qrym/InKaX6fVJ3zQTmx
aUibdhhbvbTHTxpnEtbYuAF9vE7ObsIdnajLjqxcHVTLwrBMr+SOAcTCfG+Prix73rtFere/A8F/
Yv8CU4G9b4dmnufMiKgZVPr0fx/aWujOuBvtwz4ohdvelfuejJkBXtihH1FlUcnvnMZqNHUWBBli
D2jlMPAKqfp7Tl3AbG3F+MuxFLXOPdMwxXyVzcb3HkMZwo4QJpGtyQap8AJceqUrwWe1SWdn7ZPv
sOacibEAMAdUss24z1OPUNCnRjCqYKHcZN7khwwyItLchdNdBXh3mPYjKNho+g5xqXS7Gb8F5m1x
0BJ0LCJZzSoBDlF6j7E3YGjumxZ0sGoF31GvdvEBmLeRGIZ1PpzbDUTyP6I9mnUTqwt+Rxee8jAe
nYkGFDid1AwpSdeoZAuALi8BgD55IAdSHpo2oJE6Ed5ReMba7qIlu1PrqVkccNjmUgKX1z2aG9uC
H+FXjZj5RN5av3lOR3u9Axy/PgqshCPRklHlGTfks/M3bT2vtks9StQsyraPVCLj5vmUYZVJilVv
Hp5XBMXd1kj2b8fSR1JMqmBbeQpFH6DP8siCT65eQgDSNUe2YGOkPEUgO5IHUlu9zV5BQ8wdan6t
2InITWe/MmxPPWf7oGz5apwAgchZpvbepmBzoBlUIArAjzr1Q1nmG0t9ElTrbuwWdMxAze6b/4TW
uOZ818sUdZGlGcb5Y7bjeTowRdOU1OwlpFPJopA08RMF/dMOaEdG4ZP//b0SZudhK8o+tSzVqD+u
NvMeyeQeHEu+iHZyJKlm4OTjHGWh4gPhmVLbq0FFcQtGpOjD8Zjql89lZo741oVVZV8T9IcXVpjX
oRl+PUATPZrgGyC4Cy20XnCX/jPT9cN/0wcI30c3/cIAujlDpLkTGv6BTG1Not4u/WFBVIwJbdqr
xYrAZpChYvKw+QKkpiTyUr+ycbCu+38IH0KEeoGgzH4qLOSAyVjupRgNq37e+F1os+N/hMxEjlQw
diBa/OavaKUBAvhm6E79l/4sgw1ljgq3Ta8I61QsqXheyn5r7DOG5BS2P5ITYuhb7sQcqyDRtj8r
RGqfuEnuyeC3ysaX7LUOueY/Vyzi//EMbgB1hZasGQ+HdZjU+9/Rb2T5FfeRpg8kGlo/WQtueup8
xeO97ZM7HBmAieCSPgQQHh2gFSmPPX6fHbXNia63VsAKmTe/5cX3e7x64QMSPgox28dmNEGRfbNB
7NTiv5DYk+KqmXD4SriEwhs8HgrZgFINO5AQH97wvd6kdZoACIDNxyhrq97TMfzz23xI+w/NQKoA
Jj31nKjIH7f/rASfIi7t7/TzuxuPODqccgDDBZ5gz8pSQQzEPQ+87A6AFhXCV4R9H0LAwzA2JTkE
B9ZCBkfiJ50FhvxKTkRfoKkSz3sLtc7b5ga26xHHhU7lMtpz9lcN3LnXmHrbk4hwJDuNs8HMcOtF
0sdiLXLp2Pjupdjv/PvVNGj7MmtHrhtwLKqYfn23YuZacLg/PPbzminZ3SlO53XInG5fRT1pnzLF
R7zp8CWENXCf1GMfNpaBmsPPCzZqUJ3Yfdf55S+srJa+MmbHq+QzVtJEtWUppX3B13erWscDwnh4
b4kEgHqWMHLGPikCjrGKMvmu8UcueIBr5CEOWHN/9opXdm5anNU2ReeCPOvMB2goJkLjsCtLwpht
XTGpeGIJjDsObrdkGJrDYlIkYB8Y8iiIFGdC6F2d3mcZRtp97tqz0tH954obXG+ssth2eGH7npo+
N+DmD7VXt7WPuhmGL0a+tDnDrID6+OXhQsqn09BEQyDdAyuJHb32X9vGgrZa+ogpCnryWO05K3E6
AmfUOFPhpVAGXmDzlgNdbrcl0HWxCVvBVIxe9w3wEMAYzu1oMOOQzo7+VkGIEj2O6z2o6LS+9G94
BkiFqLVSj7Z3F0uqvxtM4gL25AS7a7mAVe7fNuZpVRJI8kAH9Ry41Siz2O8NdOeb5QzFePaTBSVE
Aa1K98RY13ioJVYulma0IvgqjkvkMiGf6/pB8eEuhvDtAyG+hUt3sq/w4GAQgHqSijUFQz9HYRXz
UNyBo1K0PNLQsvqcyuGv+uGMqso5c8M82IhM+QY15vzkt0oPKLqraaOXq4nK7GMG64W6Yl8KQSXh
MQdKe0G/3OBPUzzHeV/XM1zwuP8i+CuNolJb6OL5lpI/3pc8FX73pkrjQ/Fv2jCjZs3lu66LXKfs
2ceHmhQGruokXvRHbPvmfiKgi97gsklQkAIuwVLLqPxa12V6nTEWsOoR2kkxjYs/PZQ2bCmVuAhg
cv1EzT7Vwm2phkbP2fY9VZ6VPlTyuE5cgr31rm7n7eZIZ8BIZ3YODjuH463zZU9xulvY3/H0h49u
93UueGnPFovHXKhr0n1RqPKOwgfr6AP30S8tq8t7AhzVF6MjtbJANpp/bKYDEwgQPX6lwC0KOQPu
E0y4dysoZ9uXv67HJ8NIrQ4EwVvNiNe/tfnDhqS4cu16YFXdLsHd9iCE+xVPTUhJj4KZbQDCveJc
PPNSVxdBMOBl7aDiVW0QrgsNZYrLe98elZfYiW/Jd1UdCZb74YTzTiIt6IsURf37DMYE2oXWCy4P
5qDyi6owFLWXkp1hgjA27l2P+M+3VbdeSTMlSYMLkDFJx+yEXuFcpAeut6vYe8YMMkXTfJ+z91Er
elDInNVXDIv4hz0yjuLZAcnW4nOtBlO6SfHjY5yYcbdAFB7ZiXos6aqQNZY2TjZAbSsnN0UmFLZl
uN+JhW3td1gjYwpYmh0fYLLQsnZQSwH/zFTSAkwrQ839ex+HfSxBud5SfsUFIjLgSvCIhgT9MTUt
wbXEqFtbzd229m55T3AKb8UPHfjWrOqm+3lj86OqrjF3w7MbKd1dxPV2drybKziXenBW/ZnhEcOy
nXIrcPpu1rD1hyCh/w4ml/Gm9n2qOq/qWFDuixKcpbgNwmunbLn+ur0nd1bJuJS+KHWMyFPwuKWf
jXs99CSHEk54wJ/dgtYlCogSN74dlw4QJzhHFa3rCG44hjqUMwdeNR03e9zLLlvfM//End2aDfmK
kQAiYcEpTb/y4RR6TQdPj512tWrMwWW9eo+EDn3yIF3+/hd7/0InskCxFNp+3O1q5lYsSIUPIvde
/yHg/yeT2VmgcO+SF8S33MHc1/9PBGyOFIZYKstBs0w0cctvqCJzKTisZgGOcr7OewcBmIzzy+L2
jKcQl8p6HK9k45aZktfdx5vAVUJAmmv5wNdsjDTytRuecpa+dWqRseku1d0Ogwf2T708pxf2hkJE
u24Xzc4rlmgAC+SGbp2VrtGYIWzGz1sfTdQgn15povZ68tCGg4CFxF2UdqLGYzoyNvL7G3r4CsgM
QsbYI4vjDg6on1NlaX7Wd+9GdvhL72f5TVJLI1IfA4PMeTqarWLYBMn+UmTZuoG+3nGixrtK9sOg
xzmIXq7Y4VnpGBTbny+v0nbdexOqFQOOu/Buwj133spkipVUaNoPZZ5Ks+9GRxzREIZexsXTG09n
hht0I8FZ4ue23RXsVCs1ET7W83WZbSn+BRhdHR/VFMcadQZkhltP9bhYIajIejPBuwEtLXppqO99
K3snpJR5btWGPX0ueo4dkjCVuc2O+eFSXUaZ9hE9XiigA2eqoLSxvVfBsHfK3m/28VhUg1+F7RzG
6L+Exo0MifMSjkR766/LTsYY9v01TIOugIMOHes8B9VjdfA1hLM7jFEd0fhMkAopeabC4Cy8Kj0W
94W2JC6GK8mHIEPQYCsC3+PsUeIuhN0NyT8QcE6nS5vejdiQAZTnp/oOlD8pGNdqdM10L4AKcpYS
eOiLwBZf4DnKwc5GWMgTj7Q8/J7+U4GxJCq/99T2P2eMRl8i7T31Utdw+qeyAV6DxnMYm0g5kM1B
8nhHnDn/niYxMQ819ygIsJMO+i+PespnNYqLs1nxvygcmtZfVLyCOI0arh9IwlsvdfzDl1OzMJWo
6u/Dx8QomhsnYKOYrwEDBAYd0kZmPtBKOz4MlF86tpnZvXoNoiIov9sSy2lWX+bAfbPxa/D432Fe
d7UJKSmITLmz0HKHHUxm+41WieGaFsNc2NzplW84sK5z7xRBSOca42X/Q2mQ29j2k0S1jdWXFGol
NkUuKxuUIMu2Faull5OxytWw+H+INa9fDGvoITwNI3RElrIlxwLXlaQPzHQpTbCUMlXQ3ha1YeGx
RIeL5Gqwp2wT8+Vhg3G05khSqmxbAcvAzm211eJYjBK70p5r2Mvldtc5yY1rRnsQ0JFa0/50arqe
Lq9he/HtumD4twyfJP1PY84RMTbKJbXC1ZbDF+3g0SlWsgGiSxN+1uL4EOBeYf0c48dqfSw1F3Uh
0XLHY4Uj6JiYhvpzkhvtUp+w5euaKycg1eYlG59252Af9ipuJpbOB9T3+blAwywKIMht3UCnsITE
YxTUx4ndPb1fyU2R7gyObqg1EeD1Ag020TLIR8M/gUJ393QUMzN+vaSThVwtjRDCoOcxWXWMxFok
VQepEBxSs1Abq6vxq7Gx3ofMGlVkmkL06oroKr6IxkBZvdJ0kuSnbPHydlCmc/LlJs1r/hSXkdgg
kmGHARH7lKwu1+CWI24GGHY9cQsYHB94VEw2pajfiHnfufXeKrhVoH6mGR4dGY54qvaJTCgCTrvW
1AMqlcF60QMuA5hrtPodiIPdSk2Hb5k86sl65TI7HHItXxN26vsYkzM5y0JLJHJnr0j1XlPuxFnb
9212zpSKX2C0n6not9XqnHE7azzI2RugKmikSboCn0s7vcoL0aHTdpKhryJBNjy5wMTkrtdPQ/33
C51cy82bJMpkktqEUDESLfy/z3E8L0DVOT4ODbfl/kXsIbZap2bDYbXyCc5TbvquDItttEkxkK0U
lw6w+tc1ZsU/zH893tY/y11kubnzU4lNZAm6ZU3ql7isSw0LU0AwG80c5p4QXGU8uCeBr0QhGiEj
UVDiRCgwUpoTRANkXQ92b1glTo8BQiFbBt6+Us/bLzghErAcxKDigOeeFrk2K/bgX41qdh+n3ACJ
AU+JlBbXpiBB+mKTB6VnqZigwUhH+UzdTklQmdFIcK0xQRNaDyeRYB23SZDLM4sYcgjJ/1asX1gZ
gqH+uCXaEsFT1bmMOh8jOLAHPjJvKdljHZhjYPx++wBHcN6kFGz/gqIzO5zModekxwtKP0WeTD0G
lOJT62UIVdi51dkhYazvJcpH48nftsTxyPyKZd6Nn+zKwi1mbx4iCOX9KofLD/IiJOQMPyy0gI91
tkGcZT05fh8qwr4/9Rn9HC8uYoZ7wUIpNjM5uNWpxjON/GqQteyTcFc53GdMlk62pY8ArxHKXXlu
/Kzsw5IQT0IwyLqnpCE8FGxlX2kwkMFp1NAZc3Rdou2hYWQ0bf96yR2CngffbR2CnvO1LTqXxW6U
5Q9V4bI5kXMivoyTe3gRI9FYV4Q6FlClSf61Mv6gI6cr8L4gJqTTSrWRjYshBVQEZHZOhZPzT75r
cKguDxFUrxTTOaPu8kPe/oAgA+ONXV+fWMZ8r/BzwFrTWSZRxVuim7vFMSTf3z3TxLoRwk6qpvwt
hcRLN4f42YjqZrIFpZaH1OEles+iapVOC2Xr7NdupGRi/dv8O3vEwBQftMymyS04HNx+eIaJxX95
weg4FrPvJTSjLW0Hb6foTsn5za1oiH1YNsxRw3sN5zOr7Jafhmr5UT9NEXDQU0mSpTclp/G8OJvR
FzxFuGpfQbh/HrcPi3CHwM31k6sFtVMBtFLhSKf9T1JnYXpJQn8TSykvEGng6Mc+SbEni40q0Nby
wjOOy5VLyMBzM0ykrTPZuxeEMzr1TdwqQMnew9FUtuheqc2qJSM4vFtE/Pk4rL8aZyMtye866Te3
gZ5uK9LZCGPA/oZzOfhkbnXxSciC9waOQg3obM2Xu+W5y2bxXdo/BDXiuD9obOb9Hr6OlT5hl9A9
oN39F2n3lqaIkkPSymTfAz5nBWH2gRgudd/iozxH8Ql/sM1C8hMIITRMi1HR6MDlv3K7Kldp1z5c
w2YDCl3tmChSiJ+3fhcqjEb2Mjb+0DrlyloFbPj+yAxSSjjLtLgmFHZCmh4ZYU/VX1df39YaD4aR
NtDTR3ncQKtp1XFM2C/NpJppLJcc89IJsUtytGFk/gbjnZkjSM+nPlZ73zhAavxvp3tRaEcxYS9p
Q0p/aYkO0hFiCbPP4kbBDgvE7KqnmiNnbKwSkltuwxsLwjTwcntTLaAB6YozW32sMaDyiq2Vfd7g
ZJh8i0eRILpkExsmVnPa8v6Ks6qfRWQTMtewsk6li5lQe6TLEme8cQe8bp2UPJ2hj1IYr/2eqV/Y
y3vCMsoEy0WIlwVF9aWEmgZ9Kn6QLMIBUge9y2vFUIwgUvgbnhf+NyPH954c4g/uR/2H5In+zb1M
ND69xV9wEcB0NA+w9lzzFX6xuCdrac2hMExlgowal4E+VX7RjyHxA6O8DDXXWrGYoKRAitPJrvdc
k5vtiJ8WEaUt5cmFmO2vWB1VbkP5dAtLUmW0qXhKWQM0gY/ATq4OAyorD5RDE5ab5DtKP/SOfO0m
ScagD2gQhvfe6nImoh8CnvTYhsghQTSiG6vBq2JE5lUZqLt838IbrAay3R6LrFVNwuFdDfhOijcb
lqqM8DmcZqHuOlfq5rWeW2XHr02+UPUbgFxKsscBtc2QPidE0amEMUca71Grlbf1iNPpvfJooZ0g
dxWJjDsBAXPHXbx9DGNzb5eHbCT9FlBzfwfeZ3EVhwEeaNkzB4jmWuJMD4QZv+APrGhyOmS+gv0i
LTmeCZlzFHGJ7MNV8zLJbyXP/w51CZB54nMDPqZOacJlbqRAM0owLRzMNzvoYClbdxAvpxrQ9hEV
RL27DDlNjlZqvi66XZI1lE7RdfZ9247+9umu5m1dQtvKGjvH2BKj9MAo9ZTmKch37ZcdfRE4tcP4
aMhPP0R0LkvvZh9zF1Jk0CYTkWe9DhPkqeXvRk29iS2h+3KTuHrI7qk0embEC8snmhuN2D/LaVkq
zJNBwEe5gPgB+7iY27ZP/XUcjC1AchiyyoVIV+nOXJ9d5XKmuS0QvGZfd5FnNksqr0Wc3KrTey7i
XLCCwhAiMTSl1wZAAUy3OXpxDETqfwnFZ+FKFQxdWStZXGMI0vhyCCQ0R5x8Xcj3VRMt0V0lugW0
n18OxXFLWviN1oCzIbUpSpVDJuzmHXnb6/idvQgD4s+nUvdnL1P8h0sfNlwlPHd3scVD3rVqvxTW
knNIRPQUvnAenM6uNjUryQI2wk3lrrIu7XCLquDjiMFzxYFaqfothBLdm3rcFNIQEPUhBjk8wvTI
nhw9mCcK3wFusnhLjvLYYQbpUIHw+aioFrUNb8K7XQ28XVqAnmxoKfvM2UmrcR/uLO6KUT+9SlAO
HXkWs7MAn8J+kfFYuIGpxgellcZyg8uPK7Q5apKZ1fR9HubmCaPfHOCgnDrtklzu5dClpJh+iBIl
QnA1J6q0DZ5nrsZka/DF8nL/mPmDS//RzQ3fmABUkLRx1/YY7qg8uGWaOBPjSy/je9PKThcm3xMh
9nqUhvT7tnSdMlfdmtEJLjhwbRpyOWQJNam7yRMeekVC1QSMDGgxiY+mdoh00KVdjl20hxGBVvu3
PcFxZA/EHYXOYlRekjLeSLs3tUkYXnw0Ig3IVrY7zJs7HsOKtYP2eU+2tNS+JOSKgkwW/fRPPUK0
994+l0CTfJuARN6kJsREv1fXptLru0KjlHmIFUTvJ2DWgx6viCh5rIUU9DPd9jxDr3e6mgwL6Yni
uGejtlFYkoMyiUTgtMudrl+1LuWLfVGT9E9CiIDZC/nAkLyn11NcjMc/UIqGEC1dsWa+2Id7t6Q5
3jY2+b5Et84RpabAuxoE2CG/A8HQxPIYx413id7aWAQ35G5gmBeUXdg6HpRYn3uQoWDI4nYeKZox
SdGTAIN69XQGXiaZjMqVXUN0Fq1dMqDVwDXIrM8vqv0b1HIYjJ48GqaAC8VZqWKSRwnrkI/U5US5
wd8OoZY1qbcRyFwi7u7ecOb2gb5P9iFI8tOTEZWyWN7KQI2jPhsFNwWssIYZIhpuCq7Jus3X+qts
cq68AVXfUGlL1xryw0zNR20dM49hwD9lcC2QRv9jQzV3jvlWRDMmd2PUlOoraEnoFrBpXGSgWz7+
g77UDWhVU9tH3L1QS7WAXhNFIWBEURbypq58Z8HFdjMolguFf6HznluNv4I8ZVs7msnn7RN3VoU8
oqXCYxQrEQZ3CGzgoO87Px3TcfuUZJ5F+j9WdZt0g7AoiqITqSvax1giLVyRkw15ZeMoxaIClCGK
KHkxRapuhqNWbBM7gxII7DwZp2jgopSh+N+UNUmGmr02+VPLTN4cIjoaOnFFwxYaANG2MhERAneJ
WQ02V50YEWtS5Fge7LXSxHx2WP4E3tGovDetFMZlUCDabLUDT5wsxQiR5jHj/5EaBLVJJB+zxQP8
OZVL9UXZ69szuf46tua3+uStCciWDxtv5H1+914hrlgjLcid123VDDYMnv5pOnKok+1638aPPigZ
VMJHQnkXBRWzbdJEniNlTMHJSQfKVvW0J649sjHmG2lF/L3gT6Ea4uYEsLUs8bVaCPhRvmUQ95a3
8hu4UT1tYnYmu19AuspCRUxXqiUYTantb7rhh8rZRIYsgLvPN3hSALy28eX9HaIHix5awCms0Y7R
1ItXSPV99//jqOWGzlSSwf3YlPAsV3O6Jt0FYfHp8rqEw5S2FMWMkbsUJNhIBbVUzc4CCeXnPRHQ
yYPdZeINoDRUKimDZJoIoEHhYmV+yTQyk9ViGxmcpIqspUDO/TKJoVmgnym3f3pY4LOXw0RB4pKH
t1Vp3QdxnZtn3WsC0s/l0uHeb73pl7ZlDJiTRTN59acOMzmivrdAOOTpaHAndu2xs0YeXRXNjDT6
nI/R9NU5cm5d97NO7oUwCeNt/nzyAYBtp3SWMcP97B3p+r3wwebqmg+1ccx/eV5o5xKOxLjtDXMP
cMMsOtS59ocitTinpODrpJZ6QMmddNjq4fm3SMqa3G47tNeJ8+a6dgjxETe6DPJm2458f865Vu3T
NTlSukz4jp5tLLzHBC5KXR7125IpLK1M1pBxpV5oVOiKqEwFCmDV3eJNDxYoIBrzvE/SrDjpEHX0
Bzphb9Oy4yjH3uBdwFXdIPJhJgjWld7Pi5WGa2OCNxKPENJriChYwsSk1jRG+H4wx8dpfXd/+sZv
1zrWW7lBKDyiAnDdQLbW/96YhrKDbID14LwwPIvwlIEVUfSe7TlusC8mDmU/hpF5oec7KYFj6ZTN
zimVcPp/2t1S218wyZSXUAZBs1y+5S1lYH2/yfYoluGRkAWbv+RyEaucsLX1KVdAu3fGHyBzNDQ/
xtF25lhGPVapoEM8U5QxZehDd2WfR/a5KNyUImlA00JetP0pOaw+5UpcYUy31BSYCwpY0kCIlXnp
SwBbMTwESYUT7J7/sU9xr4JRJHfwl58vVVeSpCIoqX69z47lxl7mb3ua1kO51TXgiDIJArSecSWI
BcBJSj3nNGqPOyuehXZad1P3q6rN7r8ZZLyZJuoWNPYg3Bg/FaXes/dp/9lPxabyrOOH40+gowma
jrGDCExqqg5AQuxyE9//mRogEeP+33K05KcVPnIIrv2mmZ9jRYH2U9jlfN5pgy6g05F1ctszdHfK
3h3yeOoAMPH0xgL9nvpHLEbMWxN3oLTnBHbgBy+ryozQ7wxxEXVBQFqfurVRde14J3ddDLpHbklR
/NXGSY3N6KXdgIJhoD1RK56aswZ/p9Oel+GqlE6RMnetnBohxFvEHgw0raBcjwbytOKy4Gzyhm6M
k4zvlqrrtjGEwpUQ0FztcROyiBGX5XdjkB0BNgGunNKaUcqvoG20n+NsRQRSXLW0z2O8qmclJpY2
H4PxxxlrGqNT3tFqgXdHbL1PiVOiqo8dbVkKKVbK3/3Z5DiaOz1LMju4Le07sxb3DE4kUsyhIq1o
cfXOgruAn5RsNSUkXOIG/t3cn3UPkUI09u/J04Uy5HuoQ+vf7worQEuC4thvnX1ePmcjMeJ4vj9b
YYj+L0qmNXVBsrEtfFEtmvWLUMFxsDiNhk0F3ITyaivN4n/CaZGVxVU1WVfg1zI0cpanfPEpSvwW
IZtoPc0SMdn4bDc42dSbjGU5ifQOCwQtHgf3wbBGQGR309WcywsQT6NpFQUrdjjdaKV1pIaYYVie
Z4RR+KqnkcSN7z+D9tLQck3tLNmQ4owZYYofTzGtzy5u9F2LVqedkWTLr2R2xrMwDWgbub+1XyrD
UoKDS1WYDKFfl2XwZWipqIDuSqfdv8vg2/nYoahxuSG+wPaVOF6gG6ZJRG9zOE6c5JLcc7wNuMTO
h6pzZAgRprRkzzua9QE6EktVNzUU4HeGJHML4JF1eGFl5WiWZXKIq3zzzpolw0JZVKBVLRoWOG35
WdTEliWZT1CZxo4bid4RoEVpeLKRGY8Q5D96QwYTsyLIlZiIAHN72gZkpMgTeiqGqoqST0NbpfPe
aq/Wp5C7y6QFidHJLNIa5NGDbjcI/JLBUkn94o9BLnneXMi8o2T5hupLO1QMrepPJeo0KSv9oHjZ
7LzhO14dNepTLJ7WjsE8YyJ8Cau1uGvv/uOvgxw6i0ufQ4A+TSbkfY1Xw27k/g7m3URYEsk4IEwv
tmsmfiShIRpBhy/gvs5T3KQSswSYaHmpD0zekPTz77pBC6TP907eJlDnp11HqBS3pGuiBO241L8V
dSLykC/39pN6vHKWAdcETMSerExcDQN8yHoCaLI/Yx7kf2X0knyGrLLtOP4cLjoKAt3N9oP2FRIe
NPsXEaFjBxd/wIWhnNZfxjtTGpi4fqFgi38DVZROV676+gWGCxZG52/hwhoYOnO5PpBAJfpY0sVt
u3J6tj5yNrXS8W8toqc2b6V5Op/9pocTXD8v1B6VyGpvBtskmoLBVY0o2y5RcoNIlycmTBHx+Bw0
Q6ACIySjzwMMTDbBenPqfRf9vR8n8K2gNTQ86O1FU7GN9K5rbVvWJALuzLEGhN817eiVLrccOm2U
pCQAaqnd2eoQbPAnoLoFKQK0VOUiTSXS4AoCym9hi54H+oBZFimVxAKXe8h10FP9+alHtRc89UBu
kQFEQiF5ayZiiEVrg/hgVo0xHm4KF0F6Zu2sF7S0ADlhsoVzT+OOUAwhwGfIPdvHYMgz26FJ1Z61
g1hfFxGBkmmBMYm/arDUtyINMJ8WCHQxrxf0LOlkcq7KssKLf9wtrR82zOOz3dsqu1CpOrZ55zyz
LUvl/NvO/yyzHIZTKIcEJxmzHKIlRtkv7czBSj2Z7mmfMlVqkPvAi7HOE66nwxEzWsgebuq62JVg
Xjpeye4bH0md7fMu8Crz4g4NXpPFWkhwwC5I1oV7PsUtbwHpBHQo4P0ozIRXeAHHzgCxd3SIEiAI
7zcbk12uv0PHxVxf94c8PuW0edBAXU/JghBxlHmu4WMYxtH87JPSrCV/QAr9jt86cQMDrEaAL63j
k8so15uykR1Mesg3nkOYNRCzDuEagbbT4fk4Ktx9tRUXRPYo3WNiM8wxidwTbg1uDQIb4jJkPJCQ
51i9kagiVRMN2dfos8a4dghdO3B1008B2jotmNUKZb7VuqExTvluaebI/39hlR9CN0JiuUfday6S
n6fMvyDnIXMXhK6Pji3BV8UKo3NFSNCEBwWAWrz8lliFd85vk3wOjnBjNL1sOYT5ENyXu9MBP5w9
kmt49QyQPqoj+qzSjNZE1oZ5U+EUSXozapEs2P7G+mwRqvcOeMwb6Pp5P1WjdPSTbCBh+/1Rep5q
GHtetJDAeVmKmGGd+LURoPqZckTDvH9l4S4+5barwpujUxKKYmSSlLcmTMuviUej+n32BA/mfwlD
XAVl2ny05AYMTwRaqW7mUkWQh5Eiw2XxZddM3TOHLf1E5YbQKKqjpfaYw8JhKrX5YkunFcJ/itZP
ftiwv+twzfqCj0it632cRV7lJ8tx6dwwZI4dU5xP7AIA1AlDVNkMAWdHe6fhz3Mnrz1lJI4uvNDj
7jJCw1H3b+/nayTjdYMYw9OCACupQ2LqUOcZsASDg5ZAY9LZWCWr/kC62w/FLUWgmqlUAT525QCa
r69MCoSUefbY0/ort3+AFUy7VD5ESuoGgv4m/5h6NNW1aTeSVs75E/ZRORqDhdChr63zOfm+5rR7
9FD2Ld+12q56JtO8E9h3QyoiND2/qjLVjw1vZxOootGB8Vhqhep0ZZ69KUqw6vmfwKJRVx7bgt0z
MfpBpzPjfeBbuglYStXjk0jsImBeP4bxLZREcft2B1OI438ZofdYZOWzvaxaqVMYE2ceR1I6Y2so
lN1KC0HDMP1plUV0ZdFrg+ssMd0w2AP1ELnqwhRToGu5BotmwdA58YgzFeEFblOp6oS1CXziO5ZZ
VXxCbBamo1zLxwCjH60Oh7lYvAbgDgeshtaugaBxF8K0Fu7SQ2VvfxL4IWuba/pGwMQWpIy0FS7o
uWUC8P71CGiWqv4OBCyw+oH9hEcLIts56yNvXxQFsQlqLc2Uc2Otc5sT4F4xGBKhH7wDMM3s055i
5LFPDnXDcL7ZGobA5b22qyKD+b4jpybg+KHwvgzCbqo/0zQwbVSP+ve64s3k1KrZp0CIErIpPHck
jUlKC8lVHKQ0l5PyK3DZedySQTIMZ+AuzliEvqXh8DuK90O6C4bkKkzC5gSANWZZD1upqGLtfKnq
VPzCXo332CgMM3eDHdL+XanhsfrtHwIYvx/W6JwAAfiy+xdzSJpX6OK81DVBE3qlSn8m9Zyuy7Vf
QIotY2wZp4cekxGodukla5x2rluyIi7P9Z9ASmwISaT/KnFvCc+QFYpUuUcKJFbm58w+DnfV9mw7
6E8kRHmaJLqoIpeIs7nDeJh7JmY6ntNaDKonNuVT1Sru/iTM7lhAaHKJq95OI1NODI+LUQRy7QLM
FVAopWNAYXO1fNIBnm9AyKhDGhoet+vXJFcKAyVJ5o35CBMEX5uGun5Ej62I9MzJiUu+T6VF/x2R
VDL93MeL7KwFpiLs/JQsgDPrKi4QQ+IF5OUYQwHZbolTu3db7M7qUvic59HIjgGXORzL0LM7UTEn
XzKR/BEBld8A1gB4PhGxRz+vzaKMFYLietfubcvcIqyU0lxs4799wgDXY+1f0hb/MZFxBTEstQdy
AfqdVc7YgfQVTXutnjHJIjyBTb8yaPnirDPG9QjqINY6di8YxiVRhZDA+VFfgTXWYIjXBtI8drBx
JFiL8W4HFUDv3ZYJc/60VMOUosjsuUUg4j81UMhpVhb3VzvaSgUdPID7YWZW8qPgmfISeJnGx6n7
hKkeYcYa9logJ3oQONXDiTaypfwKdFG3de5Ke+/0tbNo1Ro8fYG2qDNciPyp8oIdjw9YfwCxURCe
GcHuws776/A1MuicUDoxl+p2dQFQVf6TtkCTHvg/Am3dRXeGlZ6XX3LJj+DCB3XqAoiZ6NT/8Oak
ul/SCu5AiUZIpLzjUK1WCfk2+FPrX0FB6WT2CWsCb4JEP1058XLkYqHfxDPkBW+oAFz2NA23KQcG
3ILdL0vzCayrxC56Mzb5Y4Vx+M9sXbwhFX04m7htI7PE9VeNMb+muaNMEi/0iRd8Jq35bMTcvACk
e238CQgyXs3FhV4NYBldx8ZqxUCndoMs2k11Z1ZGC8YSx7uhFcHZ3iFOQeggr/gdB7dP+bbP6lkl
/hMgiz0D9oNhL1QnMk8vx15wmLm+y3/qg83hLZclIbLtZGkn1d1Gmdzx9Hg2dA7/KAzXWWosd3wf
oJjGpCtHUaqce3x39Cl/UQqowVTDmwjO0Vr3Xa/D63xoy6B1II4L0tfJcm2k8bitGobQmJmgSYL1
RhYLULt2X08Ww/WkY6tZ/iKGvTd2Pq9EiFIeGvaSQQpxzeuZjnpJbRiJXW2xYoNZoJkXYZDFfmu4
V9Xl8yqXZ9YeD8m5LTxp0FqtGpEQ/oa8yDxXoASjD/EX0ON4+T2GHOndRmP0OwtMDz8uCJvuClBM
9qxoiwQVQacAC3nE2AUsAvBK+ye8ZiaHcZiKJ9uhzMPOKSQ48re7epSn2giskiktyEGfCgsR4AqX
NjNBtVmvQebvakmvdkUqCuYVwpDOzgiE2gMZvE+r7+yIvyZrz+GjCq79x0J+o7V4efmwLJvbaXph
TRfUHVxYiUvfZFBsMFCaCxO27sk323LtGJZzRAUpi8cYPrz0BwG2frnFVEFqMSxJf+5cqPTn9Nr2
Jg8hexzTrI6jkVSqtAaYwtWuuRRdYq7qeqJgdaqpmm5xwYCEZ+GZ5hfx1FKJSif3vRybpDId+1Ju
aGiDybJ6W98EenmYXPnfi9YlsDVntK+sd2vR/ooO6z10c3fxTwNdb+RmK1AzNQDsd3+IedZHyIBm
IidV+9unDV9vv7Ic2z7ConTDFq18NKln0XZl5fxMdv2LrnhnqxHpMOBJoitXOVT97ZWl+eZ2HEoW
bXJ9EsnhVpqJe6vT3X2vj+Tn04d8PZOowvnauCJk7lVac9GnpsB73GdgLjx/zobS6/v8Jbz2n0Av
ixQ4e6b7ukk/oZz4VL2vEpvSl5FuSk5Z0Hirzh8Vg15smHw62IhyxBbQQ71I9peYDIcxmFqqfKzY
8gPoUl9QSwkAyH0qL2ib85SlAwNiH6K6nD8wnB63j6ZGaI9xTKS3pAwLtFCo/JTjrJ5uHtRjeuGU
GuQk3s0S2jpSPaX09tqf/he2SnNo2RVCtGCIsjsACYz9qWitQACCktoqq9lIk0n2poR0Ya08rMc0
PiXpan0dtUUsNcaDkD0nhTGROA6qzlIRCuH6kkO/qYxEbTVT4eDZQXmO3lArzvuIE8uSwyhNZPgd
IFebQD4Dgs3YwsGzIdttFGL+G9qf0IF+o9ddma4gsWd3iYosx/9Dg2V4SpeSodyZfRNOfBI7U3dA
ks5v2FpUIWQG87/BxWaaRtU/UscpT4aR7kSju3JkzbF6KA6AKr5D8HxT4jw1XzbaONtySIhLA9Wn
VphtfLAHpRgLh4un+dTr+cYeV2kEzEnuFutmJLQLOyT98Wmac18hRmNFB8eO/EtKY9n+8KHJDjvJ
lRU98NdJsBYLmy1NLKzP7VxHBDK4rnL9o0kexIDwXJrqvfZzwrz55aHXuVBJbnV1ghbA1Zibzduu
jkxkQW5x//UIKjudJB9TyXza682q/UX9lic/8AtQdPc6epasNOnkTt1X2LTcPqThI7k23JMxu1Sj
4PVk+ZIrcEAyBiXdkZRlIq9a3fRNUG0DQBUOmQSNP+YD8M0UZnU760ipYWvf71CXfsV7DqHFGK5O
vO8xNM/HlMBipeEw8rZUspQW6oxT7mefSB5Ru9hFg4l3Mpx57afuMdNr5ztq+CEVcedGH5/x03aY
+Zt7NKd/8D45zK0I58UwIMhMKZ28Ub/ZQOzUcc+IW4Y6f8qkVryiqbz/D8f3Le/j8nGI/HBjKkK3
ici5jDe/F9mf5WVECBdV8uPh04EyP27CKkaV5qfAz37TaQ1sWcNtSp6fcZI9wkQ3LmtarR5fF6hi
Vg+Awy8smvFv/3OxwyKndn6NXkDSiS7nUSipIbwty3rHC2mGaqaO+ysRJ2/Lyh6QiyeEKlXPIPlV
RTdtB7q7gd5sUpNpw7vYWGW+QhR4/GRXp0tZyZQg+KTyRXzLTkpu7/EUuzCMsQl2fDJ0SIr4f/lA
guEAIdsoMGF7pO9BNa9QTM2W+qzCt8yZTdoemm0qgiXYaYsSCxVVVA4Xzh7dKVISa1YjWHIZwWH4
3ZDTyRb7stTa9WgxKmcdv9X++Ly70GaFM7orHduoTeCpPugSLTbMqf5WDtWTtlq6l9VcwojU/iBX
62M6jCOrmV6j/6SfKseKbrA9Qg5gq3ZoqSsKRkf85fM1fkv4bD+X/Wn7fHjnIwaOwf/59abCvKmD
DbsNpuNIm7WVz7VwAx+JPBEURM0jHSkWgrlEf1xNdLdpSi11jrwEOSJhHLSnse1YysOycXaBzSAj
m4lJ/zhAo11g5eys0vkbTjp2R/LHvbIBFgOzm5xoBUBN2zbcGInXzheFraLamiB1unjZ0KFvDLoQ
C+AOoVZLx6oFxSk6dSmZsfnE0yCmeZ4Z9prW3bBAyeGvrdeF1JlyxUiUvli+x3/gxWPFsrHkSQoa
CSG8r8/IjwRpaSPoxqAI83Qy+AWqCJbkB3HfHjcS7dSnKw+d1Ja+wWa+kBMuOexySWmU4xGsGUZh
NvoJYuBWI27Rw6Z4/ZNqKKejjn6K1mmQ8Ah/CKgdWSi+0VEP4+qQAEVo41sBCPKFh1DVWQqDS+ZN
V9c27JbJkPjZKhm3jFIxV2jk3IcSDLyyEje6jV9E2d0o8nf49d6O6MIas1X4CDMCCo/2gSJjqNWo
FjVDUIyzIWW46yGzivgFwSRK45at8fn8CfIRK7KAPyWSzx7c6xTlT4YyJYVztsTxlTPLIynl8qTI
WXIQDgSj3mYrY8jQi5cyjfEvMrjoALXKEOmxnQTHd1yqAbpfZK/Gl7uoZdxedYf//oJ/+rPVvvBY
SyGy3gvgybOHJ8ETrtMVW2UGLmxStiTr15KdyhCJsf0Ed9wsIeDJ3Z7v9oIordcmbe2VIXxDm3HD
iaO/figP5OPqmDLDVZxEgP6NoThJUn+VI0jNh1+ZqsQ1N0ePDYqbDLiyt9plJ1L7Mr5WxC5Dh3So
gT1t9I2zxUFFlIq4pqh1blVCO7X0XUV2a6+mo3xhEX6u4XtQq0sLnXOFSRxkZm7XNKzNulC7+puk
2vjPdYpgoEhNEDN1kDb+ox419PeKXqd9bhucYZhU81oHiDtKz4ZWehYhS9n8aAvEBLcMrMnvEg7S
a0mn6tsHqv42JxeiMzETIm+9P/q9/+f/z5PP9ECkipmQ+IrFqw665Rdv8FMoP9pCB3DUaHX6dey8
HW1BeeQoKlaqFZSKk6l/zBVJG2ojU9nDJgU0mH2tKNG9KV7O0ais55TMyPC4GLoRCl6cjhVKvw6R
gn+CDCElsXg3BqNrhcBlxFB34sozdb6epNRVOM7pxQa4xLVywliplNVJaztTtZIw0pEg8gUZVs+X
7+4fyJPlVtFgbsT8mjAMQf8mcChH+w6w8snqpBnSoQbe4lx5S3CbLyAAnoRgqE+ocE+LPI+PMK4Y
S87FJNqb+E4f8eeL0fhrMaItFfB+621AJcuS9UtcP9Ig/NjDspXiN1XoXzTba5jTnQsMMxwA2QkE
qbuMlXYiLt8axHcwmKPLDRG8iRmYcIUqiqGQ2rj/BUKfx6bXjqjlmKQuaQzvPychD3m5QZqZGwJz
STxZN6WnRK91PoaJiZdZ27kaN6lXUM1Vbk9+PfQWNFoX+g0G+9nWFnE0/PJyOhLU0ZG2+ENUz3qG
iJdVJyGO29y1Q/NAjHQnc7y8usc22sJL/4v97ECsmdOSQPRXnJ7DMhtw8ZJspxAX0tL1UALO3PU6
0aZ8SPayxAK8RL1zS/5ysJdiiuRFcJYOX6FnLXBbDJPr7P5nmP15lTCDugXFdpO7wn7YoW9stTWR
nEHrlX20on2ng3qyV9u/zkgal72jvDWFFRhyMvTGQWlFJ8pm3tDlr8UeUIq6O0RRhBdHC+agZlpB
vW0afY+zw/NUclvBN9HaiiY2p4dj8gJYC5MbUHB0HIJgORmjLnsh65rP5wrRANJHbKFPam1qE9xR
vf4owh0OhTvCH7WC30kFzH+nxtkWBRTIH2nyv3EF8zE3wmhMLc9IEz17wVxlD7LV1Q==
`protect end_protected
