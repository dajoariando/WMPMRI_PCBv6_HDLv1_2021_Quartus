-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
yPysx4EXzslADOx74eO9R9BaXcl1S7WPKnVbsosMdZxvsPkK6xIvJlbHC7kMKREaZH4Jl3KtCuld
WVatbxMSZpfv4ne9khYECCHOOhQcFGetar+A51Qz8l6tuae0ncwrUOWV8mWY8pTGZM3jf18wRD/m
xUgu8+VjUrMb2FyxIBVNwJomCjrDLyuHOHwjDPMhFwwyTaGs8Q+WtVo6xiX7gxks1i4LQn25PVFe
UDrhnWFTP1wGeXfZc3IZuAUM1pSw+25NNMUuEG7eG3D+yheYGUX1Ua4JU96lGY6Zdgij0TEeW7Yq
0ntSTcdIyuoWv9XPZNjXcRk858+gJgJEbhwT+A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 28512)
`protect data_block
4AFO/spyqzcdDer6p52DZqq0xp4W/78OFv2+l8PRlCUocsNEY3ubWfjraey3QELQrIRH2c5cUcyS
iCaCOtUH7a6LsGRINHFi3dhMFMXBXVp3uG13nSQjlKJ8ZH1/WuU6M5lFkBAX2BOVBgGeawaUAkHW
V8SHa/bgjOSkEbCv8Wt4ctm0S7+aNyQXDM4ZqQX8Q5oaM9JH0B6nfsaBZ0khsihDudwXAvDbJpIk
kK4hZSliXhWerA2O5us4lIIMwgIGSAOi1lrUxvxDhAqTZadc8owIMR+Wz7njs+Z+XEV1o27G3hBl
tWEsmkERj6mCddg1rLAjFNmo+PhBbM/UQtn6NkVkfcV77Tk8zy1e47sShvZ0o5wDHQ7cRbJ7G+IS
YBgJ8+x6zQvFwy/v4g7txk21A7H4gU3HpzA6gli3WGaDhuY6AN+NPrkLYxkqEh5V0wRPjPn4aB6K
iHU+MVf30XviMHmz6ntdhCFpF3OMIX0c5s46MjU5qNy0fcRiujPbUckJpi/kwlh+pz7fwdQ3Fgz3
50FZIPI9CnA7kWE0R47kPgWn6wLpdbiq9aVK/ixpqN4Y/8EZyoaMymy6BnZZjHVs+v3uPGj6y+n0
RlKdwtB4JjYqT8Jqf8OfB21c03EosvSdlj839CLVtn4kSRcGkBpCD2mBfFaxHArwJQL9gAj/ggJZ
Jykxecay+gORpPhIsLHQk4a53XlwNcCLIWn4dBno6uO3y62HZaTeXSfy/02S1Tr9V9FC3uyMAB5L
bDGo14jeIKQiWYu3hNgakBYjVa5vE7mf1rmpRoU+xBAz/VvvCJQ2+j1DiKoQJ5Ri5EB3fcYuBOAL
sDfCB7fkHkoxkp5axA7660CkRtor+6jom6ldaAOGQsaS9l6zbUVl5pOu5D3X4oQHfD+U9qroFreM
ocIHZ1ZajBQKm/eRfFIEB57MLpXIa+qTluLhOnqvVf5FtYM0ymta6/Lq1tJd2alXcFI1Jpm6t5bz
6Z85RWLUI7XGWAoZnwZQ5Kq/kl4uk6owHUk4FU3fGgH7C3fXYcUelXFJSLI3QFAOGZWcllTKw40X
rI7Nnv2z+VxADIO9LinOo4tUfBvWPjR27IitXy017PGeJ1EfRzeZ7ZJ3AL4ZdJ5TYgGH4cyEtduU
t4V7tAAW+qIKXNrhBvlLvNCn4GGdnM09yXYig5m7nP0rZr/JkZfZSA7qxgNzsiuX4C6Vhyi+L+Fy
CzryaI6V/iHohHdze383FzLHHtBUBZI00HOrSbMIBPy0HK2W54hnmCyYUU5RgS/TxPsH8BTLKIGw
RqlhHMey6DP5mNuM7D0DOMyMQLJs17Bs797Yhc624dU9KoLnA62vxEjB1SZbQqyngoS+jDyfmqgZ
2qg+vohEU9QWl2pqwijdDj4bCTvtSQ6XdeQUuh9SVl8y+O8HM9WZLUHHDri8/N16xcpzsr+YOdCu
9H7Qxc6J9CZiLJxA3m9VnWB00VnLICI2ygo9TrFaqElY9GyfyxfQtfkUm+Cut7AIXUlaYnx0fbTZ
JwtQ3SjZQZNtqb4Q4SsNTQS3L5c49WKAcdvnRyGxa3i/03Q7sPf7QG081uCxOpmPe3N9VZqe8Fyv
BHFqW3M9eMBFi7S0cDmOPfdyKz0BgIh63WrcZd7mAmRQjiga+WjpK3O4iP5fN0hkSxtQDy61jwPO
UxP05FL7CwNmHRmiL+bdittpgZSyiKGXXjNSRKkwiAOSDZuDoa784hE9AidyPkYNfYUf2qAp7owm
Cmfj1qkXelidgxW427Ra2K91FlI56KMyGw1hkDr/CUD3OTLZpZvzOWH9jpv/JIKJuvKyNb8GvImV
YLc4Axt/R6zJVDo77np7eSLO1aPqXlgtllosNLTDqR6GjIMHCL4mseuL+rAIvZpRiJWhVJop8yAQ
qzJ+WQrS9xyKd1dVy1Tyn6LGYZT8QmoIWECHQx9qnf28Nixiq/w9z2JuL1Yt+Y93DAPINL9uN/97
VnOOSxeyrugFLN3cYcoGyqxgcjm/B20TYvDBAJP40Wh8Wu7vsAkff7DpIfiF2lamP1XbzHuIu8ZA
vaA1NUqwHCXntRrX5W8dDctQUb0eVDalNIu32Kk3WSIMWqjt/v2/qrT8O/auV661Fp58vrX5kOlS
w0rKzu+GDsP3+0C9muzpnQ5DANPQWz0sMOs3i72HeGBstjmVyHp2AJ5MuJyPAPXISRYLbJNsymw/
mj2DdqFxma2aW8MrbmmtC/AW85hbzUDBvuX9daiz11HyWIr5zsldnwWXGQ30hmm7DrPB2DsfIbRS
6EuMozEZvg2hPFVu/ODQrdtdCvbdtTo+i1Dud/Tt5KWcEaYYf1Y+cpdGByxMZTMnB58AWxe6CgWg
VrxaVWDmMM0PX70qZoOinC5ZT1dfUZAoYs7TATHu1t4X4vow+AKrmkISVHUdbg7WRAhGYko1VzaE
y1uRBO4G2SCCHkeF7MYQ0GsyWEx//M+jAZ3rbNgr9R4lRlCCD3+IuAAhxoUMJQ63mJuHsE/lnm87
uQRGy4rnjqwD3ji8DrI7Yzikoh8KIYlmf7hAZw7xLF9G0rc7lvBFGQKTsgcsPU/yQf4W9I+faKuQ
6zrZf1cLKhof8lqMsXj0/AHmdDsFB6PSLaYwLrWprWlmhx4HIiyCOPB5+pY7JRdbHQ7Esoj6Mt0k
47vPv4EiCw//tgFcOgv3ea2hUsOBnr9V6r9ZFzU0SaU57aXqiNEVQkF9irXtJipj5E11m0ttIHpE
nqz0ZoasEOI6L75PPvcC+hNpYEqw8i8FlpbjYUCuca5CzT5a+CNOuF/78NBaX211CS4oc3rLSztU
TbOeLu67gsuymYvDntmDYDItJ/UzEffRlQNcn0RdPJ/tcrOrAivQ+eW+c65o6BbgqDySwkv/VhbJ
0OiKGrPsFKzFOA0Nvme8Jn8bRC8UkpMuXc1ub71bAQ8AN4VU4oy6xtlG5+VXjwGvGfXT5BMyRteU
Ms4vuSUNHVGdy9kRtU6Nxnuj+mHQcqUA5foVWVgBX+29HmsoMpEU+06Ue+Z01x4nuT/AJdhPNPsi
qSjr5pnSG5tmlA9rQB3bYxOLItGB43aCXxeMMHT5iMGi1iaNFG1Q6egyhFGysSaCQLNB8hHV5q82
3hTGL4VOc6iwSTithGJtz5rVSYbeLVZkl1dCZhqzqi9fUC1l6IgORAh3sBqZt/PGUZ/Fne81/j+H
dC9m2WMGI8jQB3rozSUvpHR1IBKRZzlUU7mtiRZCDVFH7uMvL7Kjg335IPX5fOo3IZm/9sWySOX0
VWywXlODCaJ4fYVRasL3f1bY3JBH5egXBfVnKWr1W0BLtf/tvXILzIDnus1zS5o+cQFZfYD05b0q
1DYj0VTz8vi9nTnTGC3tnJuqYlqCwiTL/SXp3c5p8YJVfPNPjyfCso9ICLB69icI2orn2+uyAlm1
N7aEwh5KRCOIqKEhqkSLahcmxxReJDiF+kMDUYGAuOVWpKpobmbqp3FGluLUUepaCFFLjRnBKFFu
xr3PgYVRA6pK+QmTMNGoinCdaxnzLzwLyJzXPCtP8nm9NhIjt4oS4tL+bglE+tmjsyF9sKF0qdOF
81kCIGQy6igmvYC6qy2IeM0UY0+NWuSmgJH4tjTTM119iSsqXM3wNrfymyng6rOyChEHvaA5cyHW
yl3umec7Qg5LqED38TFEoCDd8lRxAONU/kE93/ru5e4d+j7o+4EjDJnKzDgeIpJW54OH1KBBOPmY
EUBRaZs4bg1Cxwb8DaoI8xocXNJ6Yx0KdPQscXhYJlhbYldFV8wHSdVzspiMq1zZf0FytBiDhsIw
nouf9pl/kdFxB5PLklb3mqDx6wz8eHPrv0L9q7Y08C3QNw8T+pU2M7hjsVy9TxCcanH5i2NcXPuh
o+z+gRjR9rjNn5SJFG24yjLZwUjBPxC3FNusa/7JdQxBrsHw01MbM/ZtkHfh4xWd9AnrR7Qhftu6
SdcRviBaZS+H7VwoxlYIXAtkNpfRS+7z83tThBgY1i0ftvePuLih6vTawrcm9IcRMVA3PTi8xrXW
fD77RgMXXaLsJw1b7JxlajOvbFuTO86mONakH2YGLfkthbv87hEWdQ/R4+eH/y5+/Ob3CWjjgcOY
agpz40O+9QUiao3N8w84M4S4JD9v8qyeaR92FMLg7/Sz3aKcWxj6GavwYPO8PA5/PLI1UDtOInKC
XogKqgoAaIKk0mdfsjDq66Xo6ZyQqUq3cqzv+Yk9GUoD88uksisNA6IGYsCTjYG6ECgIranMm2Hm
EFeMKvjkA3PspYNCeT2AFmU+iHn8DJDbvSZoeU/15tiaGX1K7AIgGxcVASOEltu4EcPEh7/yg660
nLlRLwJU4tTZtuuKK5Rn7su7x2Mx5p2neafjukjXAkUswkOIje1L2yBOZ/oXhD8r6aK/Mi4AgHqw
jpNMyrCYsD5GT00fEP5INwiTlAkyI0tnKP7msxziQzAkmBs7VyIhSwAX1IopgJLjAXNkD/q9ei0R
CGOsBYoE5rNvOX4VhdXqVwgrqIk1UPaCdArt20kMdeMNzTA2UoIXHMW9TpptH1cE6Vjvsvx9LeP+
cNoZxY/GKu8R5EwG1i+tdWRjpc4x1I0drjZ4ZLuF+dxSMe3Wk+VjBmCdhooCbADX2hX/U0DicnZC
qFJj9WTm8/BJw0M1ZhPi5zG4AoMCmTm+0Tcm9TfxNl285f0AQnwBH1Mpl9ehG/wJXG6O7ISNUKFh
pFbZKcvGn3tJdM3hofhgwIPeVFBhc6OaP/CpJxijSl5bXG4ag2Mm7kT4KmCwGWLFxiU9KZXa9bZ2
xEXBSU3kP2m2izPHVgPetRB2bXHqmo0u1uTbGdF1m+iGJg2gHhzg0bMy7FxgATWOou86/niAlJik
SrG252oD+89bxGa2DV8Ud6VKK5AOs0N6rBbwcepZnIuuihNgSRHuYR1UOBOAKoW5vAls1jaFtY4v
s1F2kBiq84DAz4bG52Da8A26LXYQs3bWHenUy1ADOJY5QuHf6VHuHxv5XjC/RT5fQTu7Vw83IGiT
KiQIjI1s66D4KkEWdflwR+4A+AVzD5nFOQGm7TTD1HJKNd2ZKHYTy4Ts88kbduxS+jJ+6nLtsIqu
nwmNzvq4ZSo0rquParfQe+qo+G4RpTWTcM8RxudHVkzHMubQ5LFf9CLK7kpCILbSDOTn6//bXytR
RQdBj6nZQz8Fn/tg4rnD1hgPG/cTdj3CTR+bCmtSXG6YSLzOLmcA78yHBKAFduQScxc1COzavttb
gAXeciIPQN/KeeKTDhX6PmtgTfWd81xmPdteiu8Fkhjn3ZG1A+YMocYT7xqmDivNLU7umrAaCic5
BsiTWQawktSrtF7G/tEmBkGlURY/ZPjDMuCFkiz603+/KaJiKtbpMhbLhfG25YXr3nsuwjTkESCH
Tk7gsogqklnAoj0qWo1lVKNsd9TovAdP5BucAfLHkQ7GxdC7ZR886ui8wf7SemBFmz2UzhniR5sH
4ewvxLSFjQL07iZF5VvJfXSNusrZRIfu3moM1yrMqC9v8eX01IN7wHWNpADo/+Vp1xm0bJCJdrSb
TW9gm0Wo0gHAZEdt/cYyXg9xOvBsyBkguhC89aINIR44AE0sSnXtklvcscHm4wIpod3G6jQuEtkM
b7pWbfFXRmR4jkPjYsewEVev+B8jUtCCdc6ReWbNzMwXJClHe+GCstMm89i6HxW1XnVVRLoIy6wv
Vs9Q1u7jBwkxgFWDkgJh2WRRaTW2TO6WFZZpnCCoeWkEgHHyDEljrHQPAbDnyUYqjcuXHjOFGQGm
R6aZ+wGcg0DBP1YcnVHXZLKrfc5I/uVZuQSoC64fCxUblkdvTWnHqzYngTA7zKJz8bC2APstAtjI
ivgP2C135ohOmQViThe3g5FgnYyDJ74MJzzmFMIw/gZ7Dev2B9kzKOqLs9ae5Hkp4FM/6pKfW7d+
Y+lp8bYkSSv6VyyDFsrPVJe0xcNq3tw0qSGUzHbcHcgg4A6oScueslt+JwPW6ZM0l+M5i5l3Q7ef
3Tstre4pjJyjss0uDv7TGy549UiTU/GMcdegc8CYhRJc91ccerJU1tpqo841pJpgf1EkMniC1msC
HAtIHTggihEig7r8AzRiB/igBhdgW4kxJAM6BLxFQSsjes2dGsEdXHcnl+O4L3NLfMN7qBeNGMV4
pXOGfyWrVKOlwyxlT6i18+a4tKkPhbQfbKrm9SjFxVoWB1PAEc+pyUcvN3apjlfNqXctBkgsNZa8
NRAO+bEG5hdiXhvECsPZaV3DvStzjN0LXtLlO+cc6myA2T3j1p/TiHIZJIfG04UVgdcIbuNpZLAU
tpUpttUmf7F3006a9oAflGUmliy3u7+DHcokwtBjTJy3ebf5mt6YDv86hIbxN7IVJxO8R1SKRdZp
et5yah3rBbZonV8OIhHcLFONooF9zAc7UI7o4TVxxROCgoP9/P42M/2pmjVIBk7CpSmOCFyrnk0Y
7brff+bLRRdilXhsuFd53ZU2ZdMxmD9qCCFhOSxkxmMpdRmiHBRGy2DJwMlI1kKhSr867HC+4WBE
rilqFXURn6S5GYw4BjUIDQ75cpzGbNcxTs4X05HdJ/e+FeyH1CobqbR0G24IDe66ElLOthR1N6ID
k8Xf4H5PuxmwXocskpn4OBDJgMRO1NcHfLyR8gDpEgwLNPaUeVw72SVOmyJNnohRQsKdbZFs7xtY
T0NgsLogfIGJbK0SG9HEwgpXTUIHmomvQGzq9rBz/lEOw8KcvQiYoTyMbv3nRbgUp6e0rZL6SuQu
cbPWIAPoZBOxdEfM05Jq5ccFbVezjDLEWMI+vyP8Mjqjj+Lu0hEg1JqiB/L0a6I7eC7pYqXjIPAB
JT1dpHXbOyqHqneNB0H+1ie9wKs4W9NLDOnXFy1EbwTkwIy/UvNUB0dQor7awC9NkYxrxLL98j3g
O9xFF/OCnGerTrVpEQNeSESBrjFZtW7QkarQF/NLWMb/7wzCs0dzLVW9qyPfCp9ENyCG3e6jRqMi
Jf33qv2SSX42SQaOuiHtFV32TDnJ7dPIxPOdHz/K5JXs4EFjJ0Rny/PlHSy6LU98XSJZyjLtMHyH
KkcaGYW+8vXknarhopo+teJpGZ/tdW25+jU0Bs+CwvzBooN96/FMWZieEt9GiHMhv3z4bk5MQRNO
uiJhtTUGJderTfGIviIMSuPU7Adq8s9nTZmR2kLUDOKNlGmg2Wl7myrKS0xV1+ScLxoPMN0uemHT
s4EjQGIo1G6gsJHzPiHfa8Tn3ktUf7Rmf7ZeSq3SrOcfsPOxo8AEOU36854ppDeaI13/+u4sv1Tt
LczFyFPasbMR4Lo/WKTmLgfu7HlkxBDhgXT6IiHuj4kDgaHZZgElv9NNd6JKQsbT4ZeR9zwgHy0d
S3mkvRikiVxHGLNJtiHdUhAD0TLIwZdNQ0sPr/xcW7ar4uJ+KcO5TD39SNfvegjsnoPGpYPrDwlG
T7mAgdbYPkj4j53UZqlu2JUpzMgnwU0yOLdFzGIXIgAVsfnmCwJg4yhHo+n8HLQ616Zg4X7Di4aX
6w/4AvNmxjCvUC8kaZbxqMPusRL1qHg/nTmsz3EucWfUq8+IrzGk5hWrlhmZHjo+dNW3NztQEWFX
ARA+rDj1aV9NRmsX+rWy7tchuU3p7Tcf2l1COULVmjj/qOadDadzeH8+2F1maCJal7usDLyI29O9
XMSeYqjDaXxZrjQWPyDApcgvwKBw5sw9mfVr7zkozmHAQYLHJF1u9pQPjAa+2NYiLrf3ublwQjcx
o2nfncRRPJh9IhC5LPdPBS0n0sftzBqC7DpGdUvIeiRI5oGjRajfLSjRGQBBWM9QwbD5U1AMOp+B
OyvWA1NA48U0SRbE66hWTcaUwtyP9Ii3c1p5iU0L2RbtNlr+DZ/X8uEdJu9yhNTsJ/qHHxGYaIG9
uK44mbZuCKMhw3XG3G4puVMdTocZJwJlbG1GHj8XMv0FHCUsWl0E0WxUx+uhBi7Ajd+GlykRTChD
o0bH3NWiMbNkj6CfaxXtpu5BrTLOotPEBYcCbBK6PIaOckbk1I++CSKLq1hs15PAGUAFMrzcQm1T
Tf836Z5XhonByDdEHj1Y50KbOoXFcKCriDNuGajfYS3GyxngvCLqGE7BUCqwE/raVT03RQNuyvZN
+VIjhe174H4HCYffeYSVTb/6bYbWSeoYoMvt9OMUqXMmaG9gVGIpAtQ2v+Qc19crHCPR/229VcEi
/KXe8mxSbAv6PzzG8TDbEk6Hf6/tj7Xz9smzD/0TyKLAuEeyOJQjd1v9uolzTllBTeLIjMOnmsem
idmfF4/Xx1E/bSKSCvnrYMj/OIl0HZ6Ejp7f1qJG3MCZizUaTgCCZvglEQlrO6h/+QR+qhglduOP
aXCZpUY4055ib7OLmkRlMiixjpmpeqOH5O4sD4jIqaCjC4u0c3Xk94YuMzI/9waxTNoAnmNMI69E
jKbvoP3VkoABep7AttyijRla6cT7u0/fmcjet65v8rG5TpTgCTEdj4CW/H85X8MbhqqOWOcATXZB
iUXmS8UZkqCXj0LZUdEiUg/dVDhF6a/7UgqOCPGwvQUWSN8zUczCXPONpxxpM+y+H6CZu8aibEhi
736hNBeyBH3UlL3dfH3Y9kaCk2exSR+fV6RB8SMNH5WzAzfNj1my+ZKcZKqX5l9PH1PhEv2/m0tM
7vN1CIu/sBa72WAi9gLwK5+VNcmvd6cIlPWFIQIZ046nr5/Ez+A6PosxZIm7r7cj7awmNU0R+u7R
bCMrgUBiSwAUZe6VRRPbrGsDv5SgX4mKGBwtJs8G+Tw1gT4J1O55a/parB3wwU6xKs42sk1UnmO0
fUuBrux5mYGoCOyvt6PKZbVnos6R5hwPqV9IkgodYRyCdV6J6lBdWYR2TSmvM5XFeLOe5lVKcwm4
jhP63hURqabdlbj4bOl+Qbg8MuYuD2vIlDc5QyOwV0Xxd0tH+jXtqpWStWP9IOgGiLFfxxL/ZO6b
KO++8seYAvUn8A7E2XdykU01FycJsigxEpODJqah2hKOLwcX6xg7qfWswPOT/dAhpD6bpnMmdGHr
rv0IPEL08tIHp+cE7Kcgi9wqJgkVTM3NELgZ0iYVjU0tfnkp5hpfBY7lTyG9uPlFkf68aoLW7xTT
loEKtCLwKKuRro4Zm1gcCcWmgYS8y+BpkAsx725qReJkiU6fyapIiROhZwgSNEEbHThpGN7hZygi
slvf2UTjPQe1X2FvEZWhDhOUhGXlcrEuRlV0ZL+IvjxtagcHw2dYQeMvLZr3RJAsOcgvr+v7tV+z
f2E99FMFNJ5xR7hRQqZNdHhDa1NXHcotaMIpsGMoGWqHfl9LnX4/cGLziQpolFDoxCf8BNqFCfCb
E+6jE7XehpgXYMNjreqiW1sKa8kMC10ueQAou4fGPNBZMmsApWO9RvGPT1aCaxq3jkqPzIlMkcIZ
eCAL+hv1ctmn51EAN3hCUdAiAzDewRu94JxC64+38/sH64rAEiU2DP6y5R+5GTr64dacJwjDeaT/
EXu/tV4rBB+bvQrnZkqXiIAXlD3cxvMlEM1RTtf0MOpFjdh/Iu/3PN5zEG+IXD6ONP4dIfzPA9VW
c0ZAiDzz8bRiOr9aKngDv3RhtRo0BGPLhrzduZekKtL65MF4yMhcu3UqMgLTIcLgmlWSQoJHJC5c
Di9ABulTlfjAFCH7lnpvHrIrkhE/iGFFhNZ6Uzj60fFHv8ygK5te2G3O11xjuLDPWl1YXyZ+zQyI
PmSKJNAz7dmOJvjBTEQbg/zxIu1viIxU3IhLuc2FzIyfKpxzyPr5WnWFES9OBevtur804RWsdDjA
KtsZxNwSExOfmmhxmz3FBpg+Xhxel3KlBdFcNgxM5u9MUfrNqZgGSrnjq1B8s4ax7PdfkII6QZft
N2OwwKPA5ineuN7+HfkSKyVQnPexaS397rZtqlsZNCXbF5rK7aWeY6wE89IlVyhSHQUTuoUw0Lo0
vDhh4+b1x0l/efFtqJ7Ohdl1LVH7uZflKGH8xFrdrIEtNV469qBBdwwqfvzgTcRbzk12Ws65TKaL
E0WnaBPxb7vDP8EhmKU1fis1kNCT0bRzDe1yRPxHa7QPjlc5dsU0jyvrX3MU42e82dVoOxMBQYAx
77pZmE1ZtqhCAEZTp2J20uhW6Aoi4A5WI+RJ2NtJrq/PknNHc+lMfDqF7P5bEoulvswEFRXLOarx
lKFsRxmtsSQf8vZu66A654l/9ngQEnjv4c+ukfNueadCUUF0+yq74qdGoMr+C8k8kwNxV+JfDwkQ
0PGXHnVYmgFhwKwWNpaUF/MqLJgkTQGd1PbANZ+7Y38V6uC3zOs7EGEENka4mpaoTsCbdXPFkrCs
WCbGMbZacxn+mWGALnKkBdRVAHUiYj+8cn331su1LHle+2ECBTQ2Zz1B2VitkbDhAjHT+bpg2QWQ
a1ehfw5cZr8oVaWpiZ9XaJ+sgaRvjMzgoGn3y/RZIljtzdQRxGXJlwh3S7PKwzkAFaXCv+s0biBl
BMh8k5yclHVItC0bdi1Icw0ulIEsOXcVDdOCJHfHghDJIcNOVJ05y6coCrlq9KuNfqffs2DoT7l0
/utHWtJhcztebqoI0mA+eTo7gNwXLg/1bLlLE0aCgbd0rduTaZ6gkpyFrUOT1wqJrI0bq1io+tMi
JxMq4s9YjdTp5aKQ68C+B56D2CqiNnOb0d1KmpukMdbqj1AafO8IBlDm7MJTOegI5ndBizuA6SDI
kWr5qnXdURH1wXvs1Vk5X9bAOqlbR3zfkqLta+USZOZHJ02p10UHN4s6PcIRLke5VCvgGbPL4atK
URUKw2YZrlQJqXXCvMPClZW8S6plQn4V2WgXhXRPSKb2O4zUCQfT+JxvVWxk9FUCD1kvZGlgQ39U
ivpBeMkO75Ny6j/OeW0bZKXgt+JjDk0Fsy5WgKU6SIROsZgNpZLz3xc+O7xBYq7t5O8v3KBRy/tJ
gRAENoDaiFRJmd8CjOWUVtxUFNxLBDDgKDVI9goX6R31FdVLu3Zry28yq4C9gO2SNe7uomMA0qRH
pFa3Scv401eHMVlVrUXS4sGki+Iuf3gqpzUf1wV/EWdAWjvnvHLLfGT2XmXa4GXrX6NgnKBlWM3Q
3vZi4tqsDcGCkHWEGuH9QT0gB2sJ6dGbZ24o47G3ExtJpssq5Vur7eiQFcJ2mXfcf/YsogOrH4GZ
hAxUruggMqiMJgiFtHWW6UppkwgDXdnJZ/I+YXLxKrtg6jddxkNbQ+9fdC6VwmVR1BcfAzyFYADk
xAotcwNZKX5pdQN/f/C6rt2YsXm6EaeDSugI7TxVSn9fTVxfy9AsdNcmPJ6+DhyX3A3+h3VSQtBT
OluaKmvStrETgoqSBbyRy30INtqlOLvW51e+iLyZ2L5OkYZPym/PEqiukmVDC0LqlP46X6zt1TlS
TLQXzzkhNvTnvo+VGpVVVOhS7NUGYc2bPs2PdRD6Cjec24Xa7XVtPdVWW7KyYVWlkSeU2OiyJybE
ufgxPbjPA0648QWjQZTbaWB+Wfu7sqj4npv3klr4YwRxm5i9IBG+Q3uvAQHXKYv6/BLy46TNBSZy
BuzKcxckXeL3lAojo+aErSvAMTzIT5KoCMihj3MkDmIUgF3pRaX3i31QTxJi7utYNc/NxpGjE5mu
Vj24S6kIBgHG2cIdzCv5ozRV6aG5bZQJZ/MTcWX5I5FNjTO7QeSsJmktZ7kH293R6y2LEOUjNhtT
CdLP2MEWWH8jk0hPLciOEyThATYqh3FqTlH6NWIpjzy5dWAzYNRtijkP5XnnsrJ9mtAIHNnu6sxV
HxTC0lrcrYJxHtYXcanW3V/0Pf8dK/XADSo2mwb3tYKZkBhCZ3EXqkoJcSTZP46+BR9fhePRCuu/
Zq4FC7Gtvwt3hRuhlP8A98wvaPG/vcPpl3Gu88SyrDQYkfFUjxOu97wn9GNv6eulJM5kA4YgkHgl
4g+uobzPhCtIJ+NwYj1FcW9zJ+KVlJajVb08kmudfL/tc7sbqCb6UobCRePgCfY7eDOuOJaMhQXV
kpLVXMUpH0qn7Kucz4mDyp1EROTKRoiK9C33DyjIukwt+cWxPdNJ8tUym6dBcxSxHsco8ar/45cB
jku2Rq+p1OK47L76AoN+vCE8CQh4xU9Q6p9/WG4CuYy9Bp8EudjkUuy2FLqMLC3tbfYaXPKbdNGY
ttRI9J6jBmS+Et7uk3LHFJ1IIdEN2RMn+7dqtEDhaKxDXI1IQrF6UJWOExv6e/4akBbsxNH7V1NO
FatOs9QXrDRWwc0i1GRderQ9pjtlSnFyw+FSQtH2ZRBc7wdZ+2qA0zDDVkJjJ0fFzS8JIytYbk7B
ap2UZhTBSOnY7peW7wDOqDw8QTmhvAHZMiGAEV8M+HpCCw3BM374V+OnNwZWI6h0tsb+WXAXOYNB
MtPtBAOoJt05npTTBKjHAYMzH4eCIG4Hrfe6vPUOEZ/HXz5F/Kt9aikARI0B0sIgVwdoMIYOe48F
BFfNjhGovEdTojFx8C9qEaLPZ7FNuDGeMVxkCXKvCCYNULOvqw/JmaFbBN0PpXSIS91ZjFkyEe0Z
ccHjOWtKkm4faT/plHeOS09RF4RlCjhc3EC3woz6wY+kOiP4adutPHGgPkjY0A58IDVaAIm4faTU
U0/AbqPsHaMna+xReRFl6b2c1EKq5783xNx8vAx3cv+q+he/a6AknZIfLYZ7J4+tku7WnsgMnAZG
o0mcAsvVTvvOmxjpKcbIN1uw+ngr+WMpEn5p2OY4bW6NVHu9ha3KIdSAX1aj8NspBegV5jisoWDU
1k+TU6ZdJ0WM/lMJoFRqy0riDp13xyBbQVMvTMpYt+pX7uGKWUZAsl4CGWwK9I5quhZwvvaPHIvb
Qf5Hk3NLHHB8EbsSUSbDHn71cHI/s3dif6yYLhaPM81SsSKbDfIREQCzuP7YpoKYFnAw9e4BbNUH
zu6Y4JXlop/THiIwD6V0cC33BDhivUMRJBpXXAFUnoKB7gaslqbru5lvkaP1Qyg/Y/HumTMSErfc
SHEF+TF3LN0b+WvgDlAswvK4Adrwsozuqv0GlTDDZH2wtmEu+JW2IpmRHzMJHn5nCw6CPcT3uxKi
QcUHpo//1M/FP57c2ArNYJ/UqJ9PiwTDAqX4tgsM3I50VQPMQjGVbp9uLMBOfUB7Oa0Bou2C1sTz
XRpS8G5x0WRqi7oDJj9peZlWraWAjnsI3Nwj3D0SuKswOCKGnldkf3gEmvTA8WtcQbpLPkfXYHxs
4EzVsTTp4m7y9dZyIMjrYdg4uG0jR9E37ai6AQwKU4kDF7dND/S2//jWRNTEPvKMiryggP6Yjcxx
yshKSz7qSWmUSxlblUgSY6mC/meQvgJH6c23qbA2XUXs1k0WfoVK1MM/Hqcj75sdwBcGYfXCmsPM
Yw2aZVfGqxBqCqouRetjryoSpVljy0QRHjnUCIKwpZsw3axJDPQfRRHzvoDoPW9qyvtda5Fku8yM
FqWdoL8PGAyiWf4XH4T2he/i6m/zmzurRLYmcnLXCgj2OQVM668N7ZQayLDmeorTjOOeX6S5HzH5
US9eM10nOMq72hjj8/Q6cYvb8IoACKPUmBGJJKJjrrTjA3YHCKIKwpy2QTRj93mZ3IoO9dqjne3Y
KrwGd02utqMOuE8LC7j8o5LoIIoZqIv9sASQakxlArsSoXe9otpKKq+PqYUOZItcYAEtXDZZKu0w
naBwcoCj6F+FgaGEHPGgULOBpKD5MiAW5Zt+OCgEfXVJ2FsXxIk+RexR3tjXrNZmEo1yPWiKkIAe
Qw4CiYsOW7Jv1lXq7hjt8G8j+tUMt6mDLnw1pRs3vT7wg7m2brbj0+aJfgTrEql0EtJ1WaGLlw0A
cWNl18X6yBDuPPvAa9R0cKs4HFc8cMFvwvQAt6QV0YK5K39GxFHpktfRuty1KCHSE4CBtsRmA+s6
uTgv/ML1ODzwXx2ttGs2DPqStZecRRbaBaqXHwZ7jvbBwRCdKJymLiwaHrWILay3YgFeZcGQ5cVC
wG/CkwZhbiNnC+KZxvBe2cnODFCEaIx/5woHkIrqbgaarcOc1Zf6+bj4pDTMV8cd1nrtSXJ45duM
8vghYbCOejhjg1whrNEjiMxmxZia4rywlj+AlNFq9qhDB18BlO9Q3uAW7MVdgEz6e1aBfv5/SRMd
3BDphQJ408zdZzgAJNMKvwAvTOtHxoITsaIALL+57/JtGjDtoefvmUTlLZlFZWARp1cCOAwcgzF0
J5TGfUiMBDn8rVQnsMWmMXzLR87SJDSSNffEpcmZrtsGbPoYVAfvM4wpWGqpA8uWrpfON9Z7C8yl
QHHY8uPnxYcPX7GqtaodiDHID2DKmWKeduXKQGRQ3Ab16uTwlKXHopvEcK8ajMPoLIp5BXUXHsoM
U+4HXePirdKBfMpfzZeWeFXO1XPA+Xhwsss7C+8shonVBsjP74LWGsZoB8txb30KxCeVUgv0vSdU
cWO7LCJ/v8mqfr4OE7Y+VsxuXNaUFp3Fi4xey6k1notR1nZ34Vmv1gnintcabhFV5cV55TeG24QM
jcc9S5lyZxygZVN0ZxNfhYHKn4386FWvuEpaixbKnhLLZfVNeHlPYurxZRudrpSLE0MwTlEW/g+i
3U6703285j8zi0ZpNhDOtXj5D/Gweajy64VSdRDbKsCF76+2UMOBO63Sop4h+hTZ1sxOAeMjZAU/
glxa77HG167Js7QK5KJN5u6B8mC/6bF7iEvK/RwL/3IKkUFYZApbACDZxX0ivHH75RrOmE7p9XIK
upBmTzYKbfri1RoBYlLsC3Sw1eQw9bbpWQTab+JCWQKWTLsVhGdBj6EfuRAxBSWPPLSWEo+Vk2jj
ydxOeLJ+UBmagHPvZID84x8sLJG/dTIAb6Qa+BqQ4xRU3c77PmwZ87kCSXMB6Yfi8QiePNQeIzpv
RhnW9soKZn/jqepajE72I8Fh75g1fuaXOQCSARLT1m/3Byq2wNuYhKYB1WUYwlkqbF1OPRaCuT/4
pB6jPps1Qt3S9c8jbC4ONgtFspy9bIfQ3MOKzw7nVVkSgLnnSY+o7f8FN3pTeXnL7legNMiOWbIQ
ZAEnML2fHiqs0WtBSwqwDvzwmcBYTph7XFIFAdp/uCS1TxRIsYypvv0nc2I955fSjRPSQn810ZQh
50A0pUOt67HrpmJ4ztW8iBPCDArXFIokwAGRhea0uWRok17xMWs59VfSGfGu+HcnHTAvCi4XV4bD
Fb38UTQ3Y4120CVwmJCNf7gfwI397mdtLzArCmwE5ZfQriB5hJEsq9xaxzFMxrKLp2D8jnzKMWdE
yBRzQlKa8d7Za1HCA0BTKABUm1MR4JCvymUhT4WNhdk++6QdLLMhuC6fMcnHCotx7ZMfYqb+AZYj
dthSA7v6Fec5Q8CWVCFfnrvK+XdpCc/Bgirp/tEZg6Q3O6Iquqcrxul7yvHuNQELMy1zvD0ofn1M
ahGYjAnxYDqkVhPtYPG9+TGqlb9avB0MnQtAjosXkF4cfQZwEsMVufWrR4mCXL1BthCk14W9dyxu
cZxm5Ey7N6dd8e/IwJK1NoXy6e2Ldd7KsVJR8hKaMu1huqbnjt815hAr3DuIPzQ0l1MYvAAaDu7l
TAXbaZNeftPCyUmy9i09pQxl1daTuCkbmb85lStK374mIbLLLYXtMLXmE4xWDwgUwKKROobeZE8C
JV8avXeMuZFNDYPydjgY0fEVrgjPV+BwuRwj1uF4bNVSslmfPPpByoF1Z8mjSF4JjaEegCL+J7ee
SvpLoP4AcMnHEU9vw8TUDVlPfDOHN8HdK2F6ydxRvH4ieat64eVxnX4wMS2C9rZFIytpInRd+B40
HUPbW1ywPRy5He7trXcRErWKvuY/v6P93fvOq30hb2mA7lJ1Fe9CS2DmuaUMxLsLRbp7O6R/tBmR
f9Riw5WN1WPw/jxPJlKmgOaSa3SMR6RWgFHVnL2KhvjG9Q2V78HDW7lTtwNnCp2uM7knRhfUUpGk
NAdTDK2eLLNOILqvV4LoIQBwhnCYhm4gSlFTX4puycgQyV6O9Mpmt/Lo4f+3na+RrFHZ+auw7obX
sg9Ve5GmxcMzlcgUnbYqSVLNvjYDf012BxE5w08BZlzn0autbL1UNM21QY8h4FP9s5G9qPSxBnx0
fm6pIRw59l4wohN9NIb/kTJZ9GUFX+vU9h1RRjNBGUxKMKrplU3Sfmu9Vuf2vIRlbD79GixCfi01
XAiUvjpVRoWFfaEvDt4I/F5dVzgxyx+9Ha1mNdBhrO/jIZopmUWDLwlEfol0yglNHTVZklHPb/rD
MHoIE5Q+w85/X6+57XkbeOosb+UQsnZZO3vIKFE2702Y+e23HvXs4VfeX0PJESZY0SDNAvM/aNDK
Ix+dcv0Ixv1yQ+dFuV2kbgpdxwXSmDUUGWa/jucH64/y8hsyRMXPUEBnUXZbhp/zntgNZ1B+GHuS
KYGWcqmcNrAOUH7pP9FUzT2CCEdhBVZ9zx8l0br9I+6xHEgDMYwIvCmiD/xqnYbpBi7pmqjQQLQ1
3LNMXlJvB5ldkkrojC4OTV67W66rIyc7qbcnxj1HVA7uNpQOeygnR/UAOaD/Xy578mH+t71euTNK
WHNGWS4MN/bxShbNOK9IW42j67O9SxrCM17eORd9s5nOdM9sPmO25kIunLCAGvFlcOUjGl2s9bWL
tnhraCy2jB1s7pYLt44NO0RUjP5SV7YKScd2FFfWivDzCuP5OV2MmxvhLAHSz7M3bZUu8Y8UkLb3
EX6ORJFxZiXj++MuN2PVGeniAEWCLiyiCXJDrz7Mqg0l2OJO9hayroIIPunDY3CaZ7YTSyeJlcFE
MoEShcujwKQu0Yr9OROca+WK+LEh0sVVYCfRLyl8rzYU2axEQbws+C41LaaMXwaZrT2nmfYJ7qaz
tpBaKxZDGJ9aKOEE3HIkujPOpHxA4B6RaIO8my5h/YGSXR08S/+T8OWX+vwYNvr94Dk48+zg7Wwv
vUppBQVwD9AOlSmo4ASblaTjkuFOtXNJRg4NLRaPxzQJhjz4J92jvVh8SzG3zLpZ0y7Q0pju6OOE
rVPv7V9HchFyH+/a/rkJgvqFFw4XuOE3axFTThTkkdvlx0+7CAQJXToEMskd6meipqvdvgsiUDqp
4ZVCYzH37Ni1Fa6nL7UcilOI13Y/zBmPmrRcwQqLUaKo4ovVQ8/zR298SOL/Q8Md8l2AFeZWmHTc
vwzQrhH2ZZAZcZBUjXbCo0V2ADFjixYUUmUs6MMKkkafOXdIlWT4w6zzUYx8Cdp9Jq5F/aiF5afb
aUBAAapDdt6MRz9qZmuVm1aPQ0l9EfeAkmUQ4T5OTqezMJPBU6ZPJnhC2GvDsjC2Tl3JhGCHXmNH
OOgvyIWALXtNSVdhDiY7ap9ydgTSi5Em43Bi+s6XnnGEOV3uGe0H5AkUGfAwy6+bqiO95+k67qch
X8Eg509IF18ckRwRxYlJQT4olH29YaAJvtObrYOI5XklDTk0W1EeNv9B5/VD1NIOPLdMQIrkMPdr
H8UHV+4/6mfwt6MQadNomXW2CskugfIhFkpuuD03B+9WQR05/nG4RaGys85SWjSjTMJfWCHq+ESh
X9MCuNpmmD0I0QaABCuFpUS49+v6ANKvEveh0m6UgTWKFl+ReW0dfsFJ9wXGu2sK47DR9tU9FXvQ
f0h0c8cuZErUWoY2UEgaQZLMU/2caKe428jLM5Xoyp5SiFPIa3H4PDcQeycLNbIItFBEQbAIr8C4
638z3jmgOeZm5f0yC2OWhUYLQ2AGK+iHSO547+jVhftC6Gc/OJ30mdfEubggH31N4bK1RTg9kwY+
gNhyrmLyEG4LJKNLaIxnC0c+AHOygcXR6bsabzy2YJrL3Koyd69vQ77bZUr4E6igPjBdQJ23Kcgy
NgoM9OTYf7ZjTQe/6Lc24ALSXSNxphvrYO3v3NWCAEgIwzeUiwjL8XprLJNBxxj1h62eF26476ee
odP7A7xc9gJyIAttVdqOhx8GLssyjbfbp+wXarvLS9fucFqiW7J2K0js8+IlT9BCs1hBhyC4nz6p
FxkkFCNh8MG1F+ca/9KmF/hGNG5jh56/KzrrivfoueTmiQj9/tWglQ9xTz2XLTXkRzFOlVjj/Ole
ycVD1w3Imi1BewFA4ZnUMmJWi4S8hdlqmGjwuM3nI+jfENqfaNJT+pCqT061kkgw1odT3EmK7ncJ
7pYZhf3PCt0LsinMrxJOFgSDOLPprsVGhagia8jij0ba+/hyGmqPaDj7OeiaS8N8VTFafjSMTWpw
zL8E0kDY0oN2ur9ywupwdQ15PDFGRRG9mghnwFt2j9jaCiY7ETUnT9v1H25OwwxE5/VYuFvTm3rz
zEj5MOb27Oe4GXky0sUJeFqjcIn0xBWiGCC8GOLKwKZEz+3WlDXsB4BGW+8fPdpxpKefnzdDVC/J
TG8WK5JB3BGopf/nJru4+jGS/f3RLc8g78VFm1Fya81TfnU6WGjGopUkYpC/14qyS2ywtfDEr6fZ
eIMTrhZJ7Unio6v28/esUdqi1/oY6KvBwPwZR5gXXxOHwrw5k/7nz9w/1o8hP/2BteLYjZftAHOl
KWr4/LD1ApJ8BuPFShChtv7vJs0xXcueoUrERmeoArfyNaHk2qDXaIIlRHYnFlmkPiMccd/GI9nk
3oS6Cz2lkOPvJF8BRxeJ4BRIGi0u6gZP/M5+mmUCjCKZKq2bKV9ccjOmkO9mZV/hVbN/xzDfCRBh
NggxeDWalggZ+Jqghm8EbZzeJ+iboe4VrruyAAIE4ZE3uQpJXOEWF3GMQ+wC/nI5gC527t8yNoIi
NpV1aZ/5Gk4wtG8m6TREQhPxdGB6ibD2jylaxaf2mZ9eASGlNYVg/1rRGyymduKSMLoma6LivVxX
tDGixB6jjiN4bQ587+TTxQtHUSlTLrLACdUUOhKOAAiHjD9yGOYKvjWC7Xws21HIGgWRBaDERrh3
+MOo03ggMHjdtgUTrHgkvfjb2PTZFtCkHUtlbaEJvi8DZ1IOiyI6IORyGOEOygyz9lEOJYZ7TP8V
5LfaWsRKR9qgMbl9Wmo6Kw1ce9UHw/csOhS4RiBOUPiKmSyZd4Q/J6CXmuNh4stPKVBftjzouUDa
oRWELHqyQIEu7VYySkDi44lPuBZq9pG7prVVc9RWDBMwbe162Q7apuu+/QrRgofpePOiR/Fz8r8c
gn5R6+7zb4E6VjkoZ9JPpguKdvsf2/6w7x0W4hkMNRoLYSno4rx3TqzhZcFavvxvZD6dpJ0/OCQb
cvctbkkp2A0AOJpu1YXzYjHeoWE3ISOQKJjN1z0XoeJb0+Ob/Ggd7BNObzjrvp8dA4UBaB3/e1y9
CzVdnCW4nxC64h9WB/SKuUUDEw8E16/xLXUsnbw3B5JAMVaJfdHnm1Nt7rDUkEtN9McLPBh7hbC9
ylGWmkZOHun9fNN7BzsxFpPsldLa8NunVEifHvyAavHKR0fLVOipq9+mq2EjvYMFZM/XSiaO9CcI
BBKCB5YrV0Pl1LIhorMGSEjVDAR1jdXdbsjojeZZu/QJWEau+nbFMai1CH1eU+pJHP3ZY0OwdrC+
vic2C1yri08iI6beij5Yp3OlunQhLV0GS/lVBumA9P67d0BYxZdp45hte9fjLA5BTBuIyx9yxe4q
WKpVE4wUyanaTAToP9kKz7tv0WDKudpvUObVQ+lV2q9W9ItAuO2BQPS+DzlGgg9y4w/9x/Tk9NwZ
+fr/AIxIafUlAwjL5cb82+agqO8NlN1P2LABRgduvFA10MtntVpCw98UgXIr2RLiCKKqLuaze35W
5hR4WCaVUQhdQJRURu0VIIQDCiOYGwuMtpRJkt9viStscK0oBlSpwBDJKXV5wHn3qNaKAwneyS1k
+vSKWJ4G6UuHpiWiXTnth5RmeTL/i2zbK5PD6BD9DxxLs2ONBmrUYwcqMUnmkGA27qbzRvArc9ss
f6Rsl+0HtrJyviitfDfeQrk7EmI/iIeiHeL/reg3T96BnTLLxRRQNFnb3/vtGFj5baLUbD7J87ae
IqN/6zNc9FKdNe1fHFmKMijxDNqbOXd9LA7oAVPI7lVZSBml4LAyqrqisICPzbwXxl6rb4RQj518
/77PTpoC6S6vBsamLCbH+oWSxNKKY+x+HgYr4YzP7VcHgWkNZTIscFbhtK2fDFUhXPBsPwcCAa36
1DmMRouEh80H83CNahVArFONc4Q46NxBLf1she/FoWg/fpo+toQGl1IW/zCoZxjnUUNsytKZROyW
9rDdjTjikdlRhDD5LShSmzzhAOMRYFUAM2FUsSb2p8/5xdglRKBk+Lw70zQs462FazW5Kbyp2tOT
1Fcf+8Z94t7VAGEx9FYmD/l01ZOlWrm0yAeuXtvK34CRjVioOpsef6V4KQ/iCOPgI8ATulUo8ALK
LFYvNFTCnwvUtByUCupqXKM9GrcKroIB4jek9NLrFRzKU26Uuyfm90FoMp6U62Olnv6aIE4Ax2x7
uweo92Fz7j7mVcEpcQCMIgDNyjpLLRMY3Ik5ZBQpEKvXT3DkOAwlaAJ6qXvx0H//QVZ8BuYMXk+q
oK0UBSYADsVKTEjb4ZjXDw/ZWlLEglYSK53FM9IIv+gJvQGwrvlCJcoTgSbz65WB94cRbi8zIur0
T65QWJjYXdJPdfyk54ZeWTxyMgJrlhoOMSSWAg8K5M4kKP9f6IACxAyQItr3uBd2cGDvoLUFhbxQ
wpat9gR4z3EakvlbIX32JU6X1zx+iT/d47P813X3fXtG7xzaS6MOUwBWYvuQWIiQBl7+0v6zduQ3
RSgnaUcUWIPNhjrtiHSpapAdcl9t5Nsp1hK+cI+JU9SOTWwnlY5bu6H1NaWYhaW7B494xEh2O/1U
XJAxc1lexyPKIpSZuJ+MWqqn/lzICAEDVwk6VnSOdKJzysAwkYzqsNSG2MwXmh8Mjyn3CXNBZnGB
4JcDvyztPoUUvEhECjBDdZAHWxUQ9cos95UGcFU4zqM0vgTdEn+s+xCneXFXpHgtPnZZ07UzbgdZ
Im+9bWHFYvC2wPsG8Ya/GynWQRNGXYCZVF2eVfJUyXD/cmbHx3SjaAam1OnAvkLyoimAsP1VoCLp
HnnLw5PnrO0fd3+p3BCWZEvwplVQTnJoL7Iw09qEjRIQqAR2rt63cZcHeG8mxdIvKwBTMA+3Q5R/
q5oUpVuP5mNTsNJn/8UrjrN/W22j2NXAzXmlg9icnzHL0AWB5oWx1WxYnTWsMwsxvYh4q/DHor0f
ScgPOxtcKZO5w1jGddu3v7rPc4tcqzStk0CGaHmVXqbSUSkki/KqPSb6DOLJCrnrBYe7XQDXghcu
9qIA8XknIfWNRz8ZI9gOrMokd2YzGw4tKoawY0w/9NKEPvbiZzYnCu41KR/N+WvAemQ/cgh0QKB8
a72OdQJF8mnqOo5LKQNh3LlH+5xVNvmKjtV0P6qpFda6ybsmiw9lXn38ZfiUDxrIYbqtKpmOT9/z
bJs8NZvKbRB1erUYmimVZ2CYtzlRDAGnfwyx/0J+5L14e808uxqDId7wizwIak+Sz9G4Cv+XJSoQ
Jk6ZVI0RfoCn/CxaNXS0g6CKHMNeGdxB/JPef+fIRRUPj23tL2hIhoqVEKL2MwlS1yPm7ZiUBKav
3qVxOGLe4TUA1X+GZ2TCn2YgvGI6Aatjf8KxWmUOEOOMiKXoUGUgqeOxbfNXQKUHx4/n4dcCcsP4
/t+9uKy6lYOkzFg966xeRnP71ZWZ1ZJlF9hylWBAuDY8cPWOSpjrL32YVliM1oOS2SaKXi7Aj8AB
GPRe/ENkPG0VOqX8o5yfXeCLr90s6OeXN0BaHenrpnvLysbTwTin3W5f/AUN31na/Vu1GCovJlpz
9oZbxTsfA8Sdd2QvgSzXeDubrEjQzyTWY17ZiqOpzmYKMYz00oHpM29uhvxApnGHUpcyFOBcstj/
XQvhHaqX1P7AZVLb5oygWFWuIIxODcRmZ07nkTzvoYiX0bhAZ1W/Icbn2O55JM+FTqe+s42wz9MR
ejizKYl/DH5ShVjeg5bkA50z2vwZQOIL2icTBcY/FUxTZ68Ygu50yPxVesJV254VTG+GX05wJ0fW
er712kvD+Sdn5Hy6Qse10lGb4MENe0+4F1gZTD0v6CtDao3rRM2uY7agrx87k5sgeCgnDN0iDWcu
p1s7ovkKrAdZw60xqb8GVSfhvzjOLp9teMKHonW6pbGbY/o27RW1eiI4sGfEAtGmE02+On9hpT8W
kvP55JbuKG/OYbOVY8IWxpQQnbZquZ88Dq73EZf5oH6A4+LCSD+GRyZce7lhyOvrjPV+jhGRWwJq
bJsKls2QYs691mpv02i7pI3FthMD5i5rAVhI0i6/HD5YhucOVGV/yasZlGqfNu6fnR7Zm0M8PkFI
wVfLRmZe6oSEFx7mqzWCoIvc6iocrJvxewWlji+juGq3ynCyxK/hw4WiViTKAAL01GHeSb2FxojK
DmP1GAS/gqdjkoXw2clbxhHZ7oUOcSglKYBmmA7+2sAe/+5t4JMRkbRw7lLC+1/FmNuF79XJz76V
rYxnsHuVjNkKrszyAb8DcqzmKqzumQob/LhEsicnBf+mHyYBd5qvhLMY/VfjrCRD/CPkW/Ew/LYV
/c2tu8Hc6EKp/rSGIB4dYS3v0zV0J6EDI6KW+YirjPbX2o2fOmb8X7GTSECFbmNT9bz4mVrxC4Zm
qMnoNEVfxsO/ZqwkJ6YHhjmtTEg/sTZAjtv+7PPdAvQfN8duDCp28rZvfTW1oCt/ORTTXEQosiIE
4wjxS0a1eWhrzr7c2eKUm6Lbiqfn0UYnUzz125EC6O6MA6Yu+1rsgeiqjrqiKwxq20AU+TXX8qGo
kl5ZDVpmpIkaLjo/b801rS1pCu/cBFAvZiBG7ddaKrfR99CShXBokW/XYbLX3FMBkNZQxv+8eA9e
VhS46WX6u8y/5SjL39/FTlT/xk4o9gq/etJTMKIO0Zy9wW1TPvG0wh5sNHLP9yziXtdmQ4rioY9R
C8tapodaj6FJ9KVCB81DVY3MMOYSGMtmjsUuIGCUiC8g1RfWCjp9g4c9YvNwVQY/d5QZeC/P3yvH
N+MMzKGECkOIqUD0ZGq55LBqr85vHKEuH1F0CuFC8zfGQRcuhaChselXfG5iHVTsrer7rjeZgCRO
Q/iG6pyBGHHTMw03MXj0R8n0ABD8mhilgFkLrAy31118IutVmy+DsVZmFUx/2OxVnshSE79I2BuD
w1Dj8vOX8XO7I6td4cJISOxnhKmjypJ0GWKNYMLKkTOuUAySv3/7nNrhGyKl1SOJ043Gpv2jFiRG
GA8d9ykboUNuT196IuFHVMawVweTSD47Xxawwm1Z2Csja5N3PVMHM86+kZkumOTVh4KomquSw4V/
fqm4HdFTpq+Jc6JGiqP+6QqMooL2HeFd+Kt+f9rrJHFei9w0AJ8lpp9q8LVRW4Qiw4hS8uoqLqHU
4/wp9uDUNUwiK1nQLgHjR9ItVW+Ok1kzr+oK6hQlRijD/e42q+1ia2IlP9sisb39HDQcUG1jM6gG
1mBxrgXPnalEYT96jceEJfZwHXzYuNUyMaDxyi8T6lxfEBgFHyVnRBW1jIoRYlkgcdofpqlt13GL
U65F2uRwRfCmEJ15G6zpb+EpAN/r2Mr8/ou0SfqX10m/gbaogrWmYzafnmyJrD9QTfyXFjHwwdxx
KeKGJVqhuLl9773+2WMmYuZOh2m2DVMV3/gKThoCZgTouESEjc83mFMGX4zVWEQTj1jprNZ1+rCb
hXrEXDem7U+XiMoFKck/rSSNeWE+ieZ5InWgGjN+LAIYhKq5CTzx01YrUhPqvIGGszUOqaHdVbqp
OrgAvKBB3DGU21lX4LCVVJ9LzFxOlHv0WHyEC1ilA1Y3kp+4Z1ldJMMpKwRPfwa8OfWXRAis1wgu
mV80OykNiFWBmr0pvK/W50qwZuU78cg+L9uzLRJSHSFl15PCOtrDpredzHVptPe6MJ97MJSz4lSq
VHVhwJhPoxXmqfoZRrUUbRZWVFAdGDcxACrg4zP7wDZQWKLlelqCv/MWLcYOL1Rz9UYL8ou2UJeH
6F5dLhUO6bPOttIE9b15Pp8nJ8H3DKHV1OmffGSps6q2nEerP40IRA4Z4rJsIh5J+kZdLYS6zhUw
79o7/70TCYEvx5eU2heUp/H4jKm+rxZpWLKlr73F5olyvJLfuynUgMorvgTzII5P4KgnF8mDhFhE
zRJ9HctRFYFaKe2/3TIk7rEzzXv5ijNlhDx34Zkq4+3OEvctpY8rl1fYvbutQe9LR/hUzxosm7rP
xoD4mNPYv+79o4y0jUse4UfuPBTqMhP6+4Ts3J7zqORl+TgDP2CBUuizLXbwOD3ZxBRTRxLrajTr
GSkC4ToAtoR5KRgLDKOQH5Q1VaYYMVKXiDvoBSoaO3jOaAb3WWxtBFl2C9t1GWWcDLYgr70PICff
lN7rcHAsN+ut+BKBlxBLG+qjcflidgcYHDRoXEIARGfzCYhMwLKajWOxYCyZV6CM8JSAe9FffQ6I
ADCmOvZCErv0CFMLXJh3UARQJPtYMYiBs41cKKJ6uD41pGf4577hi/FLj/CILQ3oR/TdNy5a3WE9
bsV3F6PXyJHgwq9hJrUofxQC3n8KkBNscBhaSsIynizvYHUGy1tP3kA9ZzKycpdZSTDCBSP/GZ7v
giulr0rD5Ce1Rt2gl9AD49IVR4t7iaLCwUhvJ30mpMAqt+G5iGzajw4tp7QjtHrKnYQ6UYxGWhOA
KG4jgk7O0HGGz15KDpuaLx0EAsaEb1T5iCL4nVEiszqbSFz04ZXOY+9t+ryCRb/rmRoq34axlS0I
apI8lYzl+SEXhUgoqvGS8knOhBshZ+1omOvucuzKXvDg3OPL1CpoJG2jfhfOv66uFLibqyiGsWrO
SjRVv1jFSjAI471f9Abgko4q9tdfp3vR90ZB29IEhKMe6BcfjnHr9P223X4hcjGXOk4lWia0YIZ2
LW0ywUb7721/5/VsMEfBzZ7mh1amtapXUQ9OhtfGHFdyit4TfQOvktwWfH0JCpj81sqtTSLy7LDC
jbNcS1P1a1R4czpyt7X99L1CX/SxdlPWDCcT8qxoMUSvmLvdzYvkY2yfUvXZic6Q3Fzd79kkfSM+
WTFKdKm0SA/UjTpM3I9Fcu6bClZ6aQ80Y+/vd9/fBVcTdPwpR6yDCeg4OQbtSlUwQj9xMfeCGLp8
LAOkgUZBZlUG7WercC+zcoXiuiXohYu9PE5dryvHdG+JHjMS3v09jJYJrL2HHYG0H/YHKR7JdQXq
pwNzPvuSKMGxAyTwZioDsikCCzOJPkCP1t7RtywN+HXECjz+Dn14huthKeGNqIOFHVPvb+4cVtBY
CBNNmNBnj05b6q/DwRTi1mSF388zFfw0vuKDD4ksuqyxZ1myWN4HGkGiMtLDSRAYndryo1s4G4cO
R4iQkUbQrs4scMG4yfvjDsWbl4jjLbTXxDQgUNMMA77ynIXVVz54uLQISe4Cu8LgsUdSaZ3np78P
A0iV2KE0iOWn11WwxSSGF7cfNp+cJNkxIvX98NPaTU5X2/lkCxR0R9dyNfOOEXdiPcV8dixaR4Qq
1K4OrAiBI1rcJ86oXIbPRQBOZN0Cwrfzz394zhb7L82XzTy/Q4aEdqs780MuGbWJWxOnVJ76xjt9
Phnn0SDO2lzKUO605gHM5A3fB+ietSh64/+n4OIDh8idUP6+ihsIaKtqcIDwCw6HkaIS5FQOwDZ5
Chwjcl8zVGM6OnN1KyldQDHMRYDL9U8q31S2pxwURVdmborkY5U0CQ5HL44FKmBW+gZYQrXd3fJf
Lz2CbhYJo5zBCsEz8r8Ce2ckuZulLRD4R1FExqaRH09+OgfShuyJRBzAduApYvo8/DLaOfEUjGzw
V0gLhU/fW8Hxbag7nVLIwR14AaczV89hNBuFwITtqiG2qBsWeHMSZAJbubFpCFlSJOxKeQxXVTvo
1Kpe+emfIRsHRNx0iNJhor58z3OacuNL2ikHm9Iux8lDOchi1N0wEIc4KTq4ZlvXl+ySQecgiiLq
fBmqO0GMi6qz8G76+3d06HoNdrSL5a4ImtHxMD27RI347FtsWg0ERQZj1yTxVTzn42DnYMwcqinw
XixHL0h7SCxohsQbdIM8qkax60bUMQGy0WGzOe6StEg67odmHN5GVIyMC7IiqnkclQQplzBUki7o
rgcQG/EusqGHcn5B6hfxi6ObJVfNIGG3MMBXZmWN1FyqJq7TKcBWOHqMLijaGNb4LdhvnYydi65H
Gpkj0fzndG/9s61H2EFDuI+UrZ2jkk9qp9N4bIMMg1x2dVuP/xXdNT1Q4+YhrNyxp9FD3r6BroHt
YN85h2Suukt9xTKZdOCXqU5OLMGd42PNlEmk8gCrukCKuPfYKtDYVtDu2Sjh+wkBKKXYNUSlfRPe
LS9US8/bQoUZ5601bPscbgsZpLzhv5e4CkRGModGS8FS5reUWJFTRwmQPQdfZsfIRT+AlwhWBeVb
f49H3Sx0AeN+jU29v8X1clsjXilFSqB3mgUdK9y2GjiMyzXSRTyYQYnd0uS1VO8xUxnHLCgikC6h
zEcWBt94MLfGR2J94oNvrtYleAYafU0Z0Ds1Ld/V4+FLCCQDtmD34aGAFIXtPvM8YsfGrXG7SNCV
+sNIuAi8wny6DExlyYAJ6FTC8226OaWxkeB6rzYi1IYKhzNXdGHq6EijVFUz3FvlQGHLaHXxCLhq
RaxMp1iQKy15ctMMry05YOQdtVwF00orUqcBFsQeyzrzzDExx+xDknQy3SMgV6tj8NO0Ai+oERvd
gRYg+nZJU8edGpw6XiLZN0Jyvrv2qYQXRMFUG6yFGxkKJo3z5g3nymj11jUYY/bnAEBJTlDh/bHA
e0pwcAGrfbZGN2RWQNii9KstMnKaXnZ5SQ1WIJs1/wyRi0OVUw3cfWIpEyQwWHlVZdn97kmQf3vY
GW01vFvcHXhHjxT/FYT31ygbK8kRgfKVAWn+ut61z4cfqMj4IcMlnNoX8Ch1SxlioRogCPcgEoRL
RS+F84wlnYlQFb73XY8pv5oiMgwXQdBQiwQcjcYGSWDE1QdV8fzrdCQ3FGSdvxQLo+HXGGXmqh7L
Df4mMRnmdQ7+V+pvINlOYexx+5m67kFo9VvUHRd96rCaM2abkcPhsudqZwJTofTm9n5kjaMWwWBI
JAncytFOnFhkTw+No/6xd9L5yDPQmqgZ1IAYlCXeq163DGtVftDAugwuHhJTQoK6skL2/nuxdMxj
3WKI3YRr+5IuKBf9D7RTVb0E0+qKVO7GlfG+0zZGYq+qEh5rQiJEjUT45BzhHUQgDbt02GnNmA61
4gY5wk3TNBqyE9P5J3e+rsPnAXi59I8StbZIDxD8PUNzjUhX4DTm77alQhe5lROqZbKuzh2atr4A
sOqhUgiJOPvAIVbazcsay1rGx4SeMcVFrXbFT2Hcb84BNxXryZNSekPzdIvmnRONmO6k1/+ZXiOl
T07mp7zrF4dn36OBOsdnOemi+WKSMVLafgkU0gw02X5pPKFeXEdTrvpCty8hVOlLkfUecLfI6NL0
Z78/C2WeBxBLqsfeKj7v7MBU2E/3/l70U5ElFetjiIE/fS0gJObpeox9hFuyufoKxHTuyScQL81W
skDwGRmdXd7XXGAPv+ycL5E0nuw7fePmibKI01fw4o+aGNl5wf2T1skJsajh9dfev4oMdVGMvVkc
7W0f+t5OwdY76p0MSPsd4VVeG4FpKLQcny9b8/x1OvSgS2IxVMhLrRf2bZAZX4QQIlia7Ax/gjsk
XkPZrQsUzswY6FrcAVxl/dLiqq8qJIz8vzz+WqmDLXxBb7ydNUNy2dm68TyL59f4n55S3Aq6L9E4
K6Vba6NxcyaM9mZ0L2DHNDpnHz1wReGJSqsESAZD5pRmHyK40PV+xAWpYAVkowqCbF7PliU0IuOX
kFU4k6dCXPLc5L5YYMSpIqDpPh7GD9ibU8PJNpjnHBhsB396LQVHhXWjcWTFehx23wpBaoYrTm0D
9AGyGA29if/kRb1vxBtZnA6lUnzeuGFG2WfTq7/0pbN3UrAr/fuaQolOII9oPfaDZf8wm2V1AKoT
0NiRXDBhUIj6EavlTTJi0fL56uY/mKFs26I1ZblR+lNjxZ8g6XLyVryiju+7IPzEZ9/1CtlGvFKT
Ct4x2EnoUDe0C9LN3SI3W67zG8YooHCd180Z+nRimYF9TJUvHKswKkjTwjGr6Hc6o1KEnSLsAge9
Cc69O/ay+nZiDSoCULZQjM2H2zfHWBepA3DXrC0T9oTBiQidzEMPTR2hpoqvbd916OHvnFMUq+Cl
3gTA9suq8fycT2ds7d/NlWq/XJZCrwd2GvRjjs+C8h/kLr+FBLxcE/DWWRA+ja1flwhJOJFXvh3u
YeW9bVG5Dnaie5FvSthuFBeSTd/jWsBUb1v3yT++ePgCleoE1jd8lAxa0j4PVAuyEF98avtOLZA1
NZA1X/Ntj58H7yxak6GWun291ZEESXtcuFGQoQfz4yNkz3q7c7jVDY9hTT433SHgqMCdc/vilFhq
zRoMD5aBIqbsO57BoG4Mr2IwfxbTyCqo+NJC0TdBSLtKCRPLsXemwEL7+rAEuV0uemo03e3XH0H9
xYaAo+dl+0kwoo3Hv+kp9s4Ii6wP78Oi94b2HB7R+IyyowcOu5RrQQChd+QpgEFCyqjPWUTcXYiY
mVGR/4izRJrlA6xTYupV+INUfMtQSkOy/67MNUZJm2JVwuk3QdvSGHi7yHGNengepzu0OUahVxPu
g7MHwAqM3f3Ms2JsNY3+oIhKAg44lqEZSeoX1PzKoGtXjicavRS5ne/UBO1WokPxNqSS4yg9n8VL
43NM4NbubHCntL2Q1vEdbx0qQB6b2w9SjH8Ue3vuSt2//fVeFLYNHn+VRoaGx1PNOoT82yPRojRt
jdyzQmTByClvL3VTvNxoOdvUiqxmgdqwhO4rb3aVD2YG26vF1fOMbMIdZzvc3EBR74Rr/wWA0ON3
7M70KX+zVXGD5ax2gnOKqCzUbz65T+opOfGvt5xsdzPSRWi0kwpiQWPrjwBvGKlt7YZHd4OXStWq
h4kP4ESTc3hTIE7hyN1fuSFXwCwm7KOGSeBGyPa3mpTtSKPASitDC6bRZIwqYMltC3PsPXuwKcPR
QdhQAtPjPRIwEp37dcZQ0JyPYXVAjNEW8y7P725GMkXIejTbWMTsm1sg3UIW1QEkTjiGnvPcK1eC
+DlDLi0JACln9aOd01InSXt5vAH4huDMSfaNrnmwdBPe8BTdXCFQw61cHDwlAfEDHhGjz1k11lDh
r8fGsNn1DXaOp6VrnWQZLloyFOGKhEfH/dxLOrJ3Ye1hAC+scgW5T5QjQSSFZJq9GlebAWcq5wpW
S+4oiivxaVtAfEiwBLfnSfcAMb5ZSs/mHa6c2bodOgeT3HuzA6dWv4gD9SK1W3Z+a2W9a9aRljt4
VsKwSgx0Z2yhE3x3LrpYrwDOh9KQoejBzZ6LICnAcLPrThZpRxA+5GfSrovAsyHYrJjzgVBMXsZ8
eHjVVskcnhvymSqUVuDnM6o/j+T9AxcrtEvslqw50H0Wb8bWvnZ1ozejlTHYSSu38pPqRAgTULkj
oCxTz2alIIzqgnrBkO/PLf3A4whu+pSAKFW5e1OTrAXj0wo1QI8J909b3937TuVXE+bNvbtyWQOj
Okar1aRolVE0HPaCST8iOT74Ifirwf4rNJRCi46THVziB10QMU8wtRxvMHzBsKBAO1+Wv4sdJCtG
r1vvjERMDqttW/K7+7A2osQUvMTbE1PXzpuW7GaH/ovd96A9qmr3xxP7D30S2Ka1Vf9IP1jF+oy1
vpXxK8OyzR/OCjDyyIAfvUPBC4EhNATOixkC03wLz3tBp0wMoBbrgd1WN5ANTeugDeH8+SnTTYs2
1WtbpYLRIDgft2b7heayGT8eMeIASNJ0UeZ4/6/jP+u54GDjFbnz7qqasaUSexnyWaymACR56521
YdcZCeLdV/4ZXhK+hxlzoAaNBk4LjWfxs6gSl1F1R2fRbNR3cW1n8h86leX7zn0xMc3igZwdvIfa
jZ0X5b9t8F6vryXM1lsufw/bCpwfMPbr+0EkGR7lfxkN70balQ3FOuXYPMeH9qKzLBoedCtHg38Z
7GFALixfcNdVFjybFClyjxn5nm8Cude3fgxocMg8sG+vx7p0pAiPhwk4Hodnyze6pgpSqOYKRaQg
97YUo37okGRp/qLxJLXvXYSn1HMJViueKQPDJL4jtK/4Dapa67tXuuJ8zTi7KcvUAoabvcL4g4Xf
MUAxuab6HVOyKmZxvLFKDNwpdywlgbgPQ1WCi/f2m23447K/Wj0I0PmoByUiFWSRlSr5GVLnB+9C
mN/RJyqmSBeeAN4cAo9AIUDcY6pFZCpB29ZtsXLp+UIxj2H/UDYv/O+AfS20uJ8HUBg4ic58s0t4
2jbQ5L47vfOwGrJ4K71Axw6AcsxMminVlLskXGIoszlm8cIuXVcS7Y0eO5xNZfEuAmDZEWBotPgN
U3Y/4LabnL0/MmgdOw935WAmGCJtk82YDS1AZdERiDtehkFnVcm1OQAytu+vfbRQyaRf3lx7yTD2
gJsBAWJaBOoyV3qeWxU09NJ13QMQXGb2fgHQHg0bh3n7fKwPAnOL2JB50hbd2RY1tuzgofglDpjo
ndpNDVTqJsH6HJrgji3A+sVpiRrqgrkCSH7cCIwlqMuBHs0r058qb+QQnQ3w2o36iDs/G3+QfOy+
8kWAJzD2HtI+wHk9DL9xGRL4Z+KAZ9bOk0QPBvaRATQNppeN+rmOYe62VTH1JFRZRPyFkjkbSpic
foIJSQk+R+yV8LkmVx7JkFny9p4okkPI4+hTFqPMJljkNctRTAJYrtsTZMzIovusuxDqWlZ19n97
LSi007wmhyA8kkVSPf1iJhfj4a26CTkwf2FXnOpR46HG1av+ADMCGQRn0y2++KnNLg8+cKgMeeZ0
2vvo1XvdmAdyudMd8WOWQcwMnG4VIvg8uJaSsEERT8YQ1K5RHsEXjAmpxh7fmYAhbdpn5ejZw62l
2BgkStyGnV6pjazYsUyeyUUA5IE703D8yzfzfmungnAuy5XNiN8Ab5V06WAuLq0jSKJ7u2h+UeaQ
SXR3/Dsxws0Se0IYz3rgbf9NhL8STJ3VFKu8cOak7I01ItUlp0hEkjFukEpTfbHMOazov+KlZuR4
X7L22+icXWZupOEFWwdgLVqZZnl/2dNAOlGZD9+a60MNShKkE2bmQfFcHMFY+kVRRkBoEdQT1HVe
PVCyANHTilg4QQ1yrvQWdzBEua213HWeU/iDlPQ1FvBeAOwskrbXR5sdOjiBgASGQrniDXEGYTfK
Dlnu1evq489BqTuQ5vIXiZw7ITCuFD5CwfT3L/e2pQQaAI1vbaPrpbHxBP3YTcF4joUurDwYYvRv
QjAHsue+K2z5UQb5K5bqeu7t80MlKV40duzno1GtLzlJd9H1/pxObkDCFPkFdirfe9fqXstiojb6
PsTgiqc8ZDaZ3RJR8sp5+xHvUK43bItjSAaW7gQllnBzsc/DD4WzsxVKBZepLyXRy8B/EKl/KH+m
QvcLk0bt0hESlTySMCIutQEYW/dAedC35vTfhYWozk+Fe2uaGKNh0mPyd6OJqHUAkFG+Tj0Ij4GR
sEZJ4CcoZD38RHatawSK9CW5osMjDLHiNqcclG7ikgtuus3sl9mkNZfITf3O7kbRlaU7Sqc52Gf6
GS4bGI1p78qGskFh7mrVzARtPQH5rBTsOwDg1H2S1fbSdzyEahjtKMfZGlL9jS90CDwt1HkJBlbD
3uKVsibXmvjclssYKiP3VWy7vLe1bIrEvZAhZa2NIBZV2yQxi2OThqKN75pmN/1VBo38ep/Nb8Af
BfbQs/t1+Pckc9B0EXKV0HeKZnMb5yvBmz+ePD6bNPmnGts8LliInRqvAKxv3LBMm15tUQ5s8PMY
dTXVYrrQivJWqkufdfPOcGWrSgXBIT9IxR79bojvMC/zB7nKGgcs/wfbyTLLHqDqXKuTQcHYwc9t
ULSVfWmw0ovmu5E+AET/bHypRl56K5KsO2uQvNMPjubqhpCcmG4Vfpq+H+Er0ryKjLK5Vc62Z+sh
W/9QQ6IMz6eVyjyHjoIIhq2gdqb/OF2EtZsGretNAzNGgT2dnsAYxkck5S1v/Y4oUKkh5xpFjFW7
FubR6AgiIBw2xQb2M9L3ekqJxHVe5UAIKlX9XV/wnr9+4wfg4F5cyoQpwxuWsQlR2j+fwfBGo7co
cdILtkscxmM5bhjxydpYL7jtT6ux9lhganmbKKJdBRnPy39qYOwHhExLwlhTe8bCZHONSR30nrJR
rzpOz26kTPDM5VBydTq3SlGHt0W3T+ZXGzPyG2H3mXjFIUTf0gmzi1jujDJUGj0/kdjMun2DHEhR
Nf8kVbV6qjGWu4smpFPeXCe+tDX6WGvgrsUmSnlNx+LUTSq2EGFjre3rKSwe1aJdJBpEb0zjm3Vb
43ZPv2ybAPMAiLqtKcbwzana3VlfD3CtsUcwA9dWxwgeG2uqbRsJGCWmkhTBoV+npnXTJNnhFgtV
9P5kb+ZXrvSePE1gPO2d8RZJY8kFLhFaynQ3o1LusIC2VXL+vXJFyq+QNy+f/hiyfypDJ95Ty7jT
GPTfq27gYLytiVfsLY6juYDD+96GOFidD7X9uQIR3aM2u8HSYK/lzqJM5JOkD4Rk1jR6zCZxjTNY
aH7JM3jzACjkUfVExyck7TRoK3nLyEPQmzA3Jk1CAQ91MWyPEc1xsdfFmzmVMo5WkquujM6w4+Xa
SFYRzlWcvzmDhdVZeYQGIQsW89UpMlKFylBOcweAQThm52HQ7gNpjNmK5z8G22trwsQi94+NKi70
LSvrGkRJKY0v5l82NUOwLh798OpFgTSSYvz13xtH23QKxbKI3XSYZHSSm7Ggn8GdJPAGzEYGd/9N
xqJ1miuUxaBrdOxxcSPYx0CUsL/3su0WTh5s1SdPbB8V8hplwpCNB0e4x4sCu1aqpIUGXqpR9OxJ
Fh8ISIe9aAjOSqjrRfJx2pDCpP1hiia1I9M14xW8O1QdULlRfa9bdwhfphNJoYkpTn1XpBm20okz
QOXwz6MRASWrT19HMg8s1TsualVe1i+QB3CkiAxCVTa0eVdmrT7TmsaFqSXeNZKXpUz8WNeS04yL
eSFon6qtt7+oGJEAPISscJiIVWuN/UrA6a5gxhxgNQ3+qOUdBcHrc7MfBmd5lqlXaAsalwm/LcvN
+AExJRz0XGb19rLMnEFYjeYl+jbVqFeJHTBU80Cqim70MLw5veJISkwS315zKfrwTD0eiBFZa81o
7vx55GFgb9MGrwdpAFW8wrjqM7g+MJlJLda5tWDp/wq9wDuTiBwCWTswNKGQz3IWHpkPPOOEFBeY
t9HoZSbx4WJam7ig5r8qaNAuaHVZuHo+xRPu1prjkKfOHnmjDlaIhtFhrW0OEfYP79RzZXRYxoUV
K/+r27dYgJyIolwHMWGUhXkZ8NXr43iur0cp5kOJoHuWr3okS9sQ9K1BsiprlL6iJ/SD08Phut++
u+k2Q+kEZ7rBrRg/ZHc+8DZ/QUSld3l1SRt4s1RYLae6b2lgwz3h0uobFcAnfwOrhei0OJ5FYnmG
YOBdzVZuamLVoBT0B3P0g34vRWF9NVGDZov9TWCS+nsKutxqXOahSpKUr5d1UmcmUfg8tOe3EzVy
JTkYuw8CNHNANFFUZp194rSYb2sNX+hsESU36+JLXM/hHyls+MxzeT8kEalAgZbnVvOnn3R8lebl
kkzBP+unh6qk/F3aNr0AWkC0apLdbGWfLSIiEyEuUKn44xdnpOUxb/MXjF3nNXpQL0A3cXIaoxUX
DJ4Kte/LettqX2U7VsbXQYhOHBEvu4R+4pGdGPkC+QbZDSfU45Z3fvgEhzmRLMFrOWGVFo69+3Ff
jDadFro6tJPRvdAQZfIkUNIq9pDOzp84Ihk+W5WoddH+rTzVrvN89tfvi4XTa8hh7KQzJXTCYZdm
kUYnolzkeWzvvXIttpn7YNmiUhH8q/mtzWkqUxBkT/D6rumll43JzAdP98eUBX5We7+oXdhLyoYC
jKVbGzwUW+LGNt84zoOhZvNx0xTPrVKE653p9KCkWBlfyr1CeCm/+dKVTRjTtQolKgCn+gPgMHBp
MX9nvcOZkebjJ8jlaENZC4n53eRgVOI/CB4p5Km1XjvAa9PLvqCVJMKmgZB6JH/fNTgodxlbEdAW
kgDXBSP+pB5fL20lnN3T4GJPbjRf5Tq2CGye8R4bl5zulU26KPgvj0xDKEzX0ZKqiUh2eeAW5XhU
fv7+UEPmQVcrlRTEXk9BilDDpwX0dHRo+jitV2TI1H/PmuaKH7TZgZG5E7MKOmIPBixbe1mh4P8m
pkI6sDuaT+qZm7EJUu2JKu26+5sQb2hEd+sWvuRiF/A4d4t4A0ghphO2m42fdjT6mVAftttq96nD
slZmmJpAFTbh9M8BaliwAjDFN050RjUJl4JBDac3F344ZrHO3AMnnA4MdeQZ55COywEqHv+vUKY3
/CsWG+p0YpCL9u5JAduQgDpYrwG/neIdrPlrjiOjx2WnVvcyJuu8TLNPjfYVdxjut/LN1ZYgFENp
Y91Mj8J5rLFjLK4m0EqNizt5Ln+mDn8XNgs8/Vr4o3GGe0byXoT9poPSIFNyI2dzFWeahO6+B8Br
fl7wERHsMPIdTL4PCPvvqKYoczIc2nYkrrxDqzB+oUECQ5rEDQ71Uz4MsYsT491z8IML7U3ErLRs
8ELZqUk/cOSTZZT7JahdW8YJZEMVvHCuIEX3er8TgvcZfVa1+HVwrKWl14odobO2NQYvxucHwu5s
iUkplJadtVW353nzz6kHdQKCQYFxEgbJDfqtGzm0jF7/LHRo2ghkAsOyYQkWGMYGkkF3C0kqYwfV
4M5zSWeTCYo4j5FYR2A1LU6TC8JKiQboUCRbXj2Ou3SFqEmHq5kSjdv9SQtlFSy6+zqTPu6yVSnT
MO/bm/q3h9twUYMv3+K1mbWlRveejY4mM6hZuvThph3Bv2/nU+mDf13dbNZ6WhJRd/nWwJ1wQ3NI
rVqZuXxEUTManKk4EbV99dEGRSKYhpdl6FHiEAKlPIGVrZIGllKSY6wuhWMBnlrLU3tVC3481+RM
2v8t8aqW822kbPsNQ6CUMxXDj0xDfMWcIt328WJZbstySr2DFsnR6wupoRsGEgkrQKYJwKPviIGG
tUQxBf0657MAlZyE+FHbD5hhANYfgA7GhV5JX9fx6YGqJnMENy+HOZBRyct9jUtHJA35lzeGPn29
vVm/D49BKEW6crdOvyhBYyeBkC5YmChrqCMW94pK9RjuRyT0oSZWQd7xVPOvGvGPTg/5nB8dJI47
MNmIDtIR3chSw6X/m8mn+hy7yAIfVtXNhKBGMtQx/5Osgoj7jsROy0lhLHFqim/kp/HIcYTTzqoi
Sk0fgmXj5b2jcYuHaUagmdF9dUz4i/yjhCF5nwR6W9nPqH/SpeTnj0f2UiKiS2b6MFlMVsa+ZJHj
3WLo1nNXZ5YRyEmz2TtJYgXPBLwGg+sWUDvDRRWNkQsuUa0OeROCOMO7VQ+PPaEF0eyCVb+scXIi
10AGtGilAfNXKNAJ94Mx88XrTvSFsuEMDiuX8X6iWGlwNI8L0Tnju2klAAG3rFw6DlSurPIwUeCT
+Fwdlmq4OJGKe3DWO78HHdzN0SCH5MNKJrD24JwoegQ19iSKOBWbFPWQLlVrrVfX6VD2ztOnza8t
bZl7VnbtI3cl+4YeXgBsvDKoVhEYdw7aOxDdjZCgSCUf296raPc6JmfSVHvAGoJTFBrMsFawaC+t
k8Z+f51Hhqzn8jf43odul8L8u+/UbH/SxnwmNZWrTkE4KkQX4j8OcfKeXQFzdnZm3ibpDZDmIH9v
YhtD9y9JcU9DrOBBU/a1o9Bfkl2oYTSXMeSPQwaHLBzfPP2K50w7m+QszcfFA8xGY7Doh7Rq3L1/
pAD0AvoeXzYOjKESzhm2no2vkJd1SOTW85DeGx2XbC90GvA6itzYb/u9x4iWFJroScVfSmVz9huL
o4AdVh6pUi8r+C2ySa9DGhtMeKEl/et2HyBy2ErPG9UbCfUlkQXa3aaOCb9IFbPyOBnENcQBfBC+
J6aH8ib7CwObnIJcgV3vrAuymrAXjLAWFLVG4y+Wq06SLGJ2IjB8w7R5GWHHru8NHbOaWuzlLK5n
/ALjn3e7cYJcWzLiJxBsWShX32G/zYgbge8y/Zwzua6MubChh55BoaSgIK4zWRuvTGBYIwLSjhxw
8V+9Ang29JowjhmNX/2tfrI2OOVRqOOrhVBoeF0KHFm/MrIX+//C5KQYgi1tXiBg3TWD+PlwdX4G
b4CqC2KFzFxnuYIpgjbMhEzVfx02+mL73+HtnKjZNRq24aNYxWV4KybkxX2Tkd8qKHn3jhSfFlmV
txufw0E0MwmB0HRbkwEXRWiXaVghwvitxergVEmqh1R+3J2a3coVBzcM2AQ0kuWEmpw+KDBJjBYc
uAtyHS2pvuivcSYzxbWZF4GCPp2D+Y7VXg68QFqqsxGzs/JvmzNx0Uk6dBUc75FNDrLmW2BEY+i6
jsn4/3bSwfYDFdPA9rNLN2ZxrthAJ29BCeKV8mCRrT3OhCsbsYUy4J7Q3D/t9MRwkdA9bbDAeyBI
KZXsZQMFA4NbLF2nLYY77eZY0af9MWgvhhEkaSfCAYXCdRSmlIqj+pJ92Dqfd976et/8X6RELpvZ
fy7oEkCPUTfoqfaK0k++oUr7RifQwHwa72dRAv0E3YX/K6LRthExyyqvr4Yy6jvaC+tPLIw3DDPf
7+WwkZQP0OHPL7i9W9jNS2trY2OtE4BnEkpJsfCdjPCWaCbO1aez4x3eX48dcbIQq3T3ZUDJlSdL
ZCETDqfHbUKWDLQ3+f3ULFsjvsQeTVU6A5/tBV7GMK1DHAAJNfSuqX67jBo0KKHBeixsfnvbgZbK
japqEM+VtRGewb9NlB74tdJitt1OerwfFA5V3k08wQ3Ll5fbdhiWFKevjg9KCPfrJXa7RCPQ2AbW
qRUgRR5Q7nQ1AYO6xLKRCHJ1i0TlCSSG6tfNBWcxhtxwUZHwPHB9mBQoJIicrvEmc3osXS2a1xbI
GIaOJOZ0fSJNU7ydcOUSFas4lKXdYoHelTWVDArcuiRCfLzzbYsJ64xOH/aWwLqYL7VCWMY4JCcb
CaoYux+PzFD7qRTljGcb+I5uMvy09PWuitcHKs/ZXCs8L/B1TSQslR546T9U6hlqsA6gl2zynrkk
KrgiZ5HNgjZkxEaiakWBjwYjwgie9g5KM9lN5IdTVdV45qI6Bqebd0vuu1c/e84n0hXlJx81gZ7S
XwV8qhVIGG7iZGPlWQF52CofRyx4/CQppBr5v2hZjXFl5IJIONJW43JjslDoSYb5h1O1A0LI7CT3
kYvcxwacfB6UV1pvuch7xE+yUbwsi7kFLXQx8OB8D7/7D3nJKY/OveS1QcZNpXDgvn/QOW5dOaVe
+NeMXfiMc2ShSFXJQdmoTz+1jYuSdpimJX8yycsVOvDQyUVJjLNWeKvzlMmlbL3nsQIP8fuGnZ53
3ezT6W1pJbBWvBsG81VsJ8RPwh/f1q1c0rU0olAgKubYwrgamUXZbiGiSZwgIKvB/RYpJmArCZO4
Lwfnyk7lq5qaFEJ8Lfp2bPlK8JHHrWzHUbulHwcYxxzReA3YtEXjXr4vL4grMTYGKVMkBBL0EF+a
4x4YtAjaFzGd2CmABGJ0OwCfQ0P0VsqE3lFQH3uoFQQjuKOSnkM5QqQt9di84eTBx7Dli3odFsJ+
au2MBH9ooNeM0jLEoZJp5C2eBKmOC3TH2I7p/Bsw75Guh1v4RON5qgaOtH2Jgn2igmfhrs3qVGNF
853MoPhTRbFu41r8AG5m0owicmAmrIPh8TG5RElHgC6MPvwsx4VaDyaTM7mMPRGSVi4V3J5tvp6K
AayoD4DdltME3xz5D5+/aGIqJpaUeEH4UBTbfgkbO7+X7Sa59aqozo19xSNkoglxaaHshwxHwdvZ
VUkQmpD7Hs8l94mn
`protect end_protected
