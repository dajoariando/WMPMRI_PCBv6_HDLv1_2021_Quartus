// fft_fifo.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module fft_fifo (
		input  wire [13:0] fft_fifo_in_data,               //            fft_fifo_in.data
		input  wire        fft_fifo_in_valid,              //                       .valid
		output wire        fft_fifo_in_ready,              //                       .ready
		input  wire        fft_fifo_in_startofpacket,      //                       .startofpacket
		input  wire        fft_fifo_in_endofpacket,        //                       .endofpacket
		input  wire        fft_fifo_in_clk_clk,            //        fft_fifo_in_clk.clk
		input  wire        fft_fifo_in_clk_reset_reset_n,  //  fft_fifo_in_clk_reset.reset_n
		output wire [13:0] fft_fifo_out_data,              //           fft_fifo_out.data
		output wire        fft_fifo_out_valid,             //                       .valid
		input  wire        fft_fifo_out_ready,             //                       .ready
		output wire        fft_fifo_out_startofpacket,     //                       .startofpacket
		output wire        fft_fifo_out_endofpacket,       //                       .endofpacket
		input  wire        fft_fifo_out_clk_clk,           //       fft_fifo_out_clk.clk
		input  wire        fft_fifo_out_clk_reset_reset_n  // fft_fifo_out_clk_reset.reset_n
	);

	altera_avalon_dc_fifo #(
		.SYMBOLS_PER_BEAT   (1),
		.BITS_PER_SYMBOL    (14),
		.FIFO_DEPTH         (1024),
		.CHANNEL_WIDTH      (0),
		.ERROR_WIDTH        (0),
		.USE_PACKETS        (1),
		.USE_IN_FILL_LEVEL  (0),
		.USE_OUT_FILL_LEVEL (0),
		.WR_SYNC_DEPTH      (3),
		.RD_SYNC_DEPTH      (3)
	) fft_fifo (
		.in_clk            (fft_fifo_in_clk_clk),                  //        in_clk.clk
		.in_reset_n        (fft_fifo_in_clk_reset_reset_n),        //  in_clk_reset.reset_n
		.out_clk           (fft_fifo_out_clk_clk),                 //       out_clk.clk
		.out_reset_n       (fft_fifo_out_clk_reset_reset_n),       // out_clk_reset.reset_n
		.in_data           (fft_fifo_in_data),                     //            in.data
		.in_valid          (fft_fifo_in_valid),                    //              .valid
		.in_ready          (fft_fifo_in_ready),                    //              .ready
		.in_startofpacket  (fft_fifo_in_startofpacket),            //              .startofpacket
		.in_endofpacket    (fft_fifo_in_endofpacket),              //              .endofpacket
		.out_data          (fft_fifo_out_data),                    //           out.data
		.out_valid         (fft_fifo_out_valid),                   //              .valid
		.out_ready         (fft_fifo_out_ready),                   //              .ready
		.out_startofpacket (fft_fifo_out_startofpacket),           //              .startofpacket
		.out_endofpacket   (fft_fifo_out_endofpacket),             //              .endofpacket
		.in_csr_address    (1'b0),                                 //   (terminated)
		.in_csr_read       (1'b0),                                 //   (terminated)
		.in_csr_write      (1'b0),                                 //   (terminated)
		.in_csr_readdata   (),                                     //   (terminated)
		.in_csr_writedata  (32'b00000000000000000000000000000000), //   (terminated)
		.out_csr_address   (1'b0),                                 //   (terminated)
		.out_csr_read      (1'b0),                                 //   (terminated)
		.out_csr_write     (1'b0),                                 //   (terminated)
		.out_csr_readdata  (),                                     //   (terminated)
		.out_csr_writedata (32'b00000000000000000000000000000000), //   (terminated)
		.in_empty          (1'b0),                                 //   (terminated)
		.out_empty         (),                                     //   (terminated)
		.in_error          (1'b0),                                 //   (terminated)
		.out_error         (),                                     //   (terminated)
		.in_channel        (1'b0),                                 //   (terminated)
		.out_channel       (),                                     //   (terminated)
		.space_avail_data  ()                                      //   (terminated)
	);

endmodule
