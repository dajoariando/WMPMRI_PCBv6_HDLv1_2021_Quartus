-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
c6Q7NPnIhtFPgavpWrpdrS/YlqwMXVO+wixOnGFecQbO/1GiFqc4YmmAIkETjmQHmOM61IW3b6WX
LW7Rv0qmjBCI36afc+xYJ7PnTGc7MUFQ6ve7+LUmd+0p5uLK3T8YKzODlu4N8cJD0itIVqwPqNiZ
nTB6B+mPXBarwm5CQHM/Z72hRV2+diOdBaagOAuzbXA//CfWwomgFWpcpMzs8ri71UYS7mxwnuDj
uYS9/vA9JFzuDBPMJ9S8i8W9TAbS+UbUB9UZTJP3SH04lPTS+UYwTTWDzmyXIAW3w7vbLp4VGQ/s
DFQ3sgummZYkSo9oI4PCeQfrVPWJ0MrMLhAyyw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3328)
`protect data_block
Lf8wNVZyXtG4Oy5UOzkLz+aFW+MoqtpXgnbJvLCiwf9/6u88AufFo8lna5IbY5D8wXR4uLu3i9Yg
jC28DhTBnVjslYM4rZHE2TS9G4WLUoPErksmViivoZU/Eg2NkNCXYHsSIfF4RhZC84vVFLGNrahP
cTa8bTDUeFdd6oe14Mjcj8itx9p0Gkcxj+OOy5E4mSLTP1FOfTRuYStp2HSaqP/ocrAMuHui0PnM
acIep/kQCYRLM+mtnJ9bQFFRyIj/wM1AWGVwogrhg79YLIihsnzzlrZ6iANAfzFNT0FPf5q4lNts
cgb+D79FPU6xnFn6lkF+JKAkTaYKAgYiWZty6zjIORteDKdsilnsOtEuCf75NElkWJE2KzzqSU1r
owy3gg1451M2rSo3JiDJ/puljwQIlm1JrXrJVlVbEJxSIHyTVUEBRUqmnbhvEYAvLg5NCvTnj8mc
0YXmTvviWrDKf7SGfz/aPD72XXY4CYuZ/25XzOTpWJE+sR4AZUuc807ANy/uAoW/qqOc5eX/w2lV
/xzwu9m4p2ylwDBLLZBLJfXy1iW1pO+eilQ0J+8qtw75ml+uMV43tqRecHTC+ptbxcXNmH9pyLX8
l14LztmdAotddDOJ2rZehidnCxMX+raUoU04zkWUGivTjeoRA2iU76Iqqz46d5ZP2ZzaLmJwnvEB
jRCsJG5eDilk913ogoWPz8NbY7/tKhpZOwbDd4V0CspkJvtQGtkMubgBqzs7LM+6KU229STwYdDw
Ifzs1Wxws0HRzzck/IyeQonnRNFrArw2Z2yDeGR9D2dlj6s3+5nub6YMLXf0VGr+nBbXRgHIUHUU
T5gh/ec3q9/oK8pU60lhJfWffLWPmuMb9vg+QjU3Xbn61Pwj/UySnHa6PQO7mxRoDoma6vc3B8lR
CZYBe61Ao3PcL39uHCciwaRAOXiZFX00yVtMvs9/SQaB1tr99DiVJmH5/LIxrRuNFxvx/cVOTAJY
+u2jTl9Z+8YK7OwQ0hmDfoAmOVDcMCFBZauIMjbNrkH+KmeGZqugkQR8IcY8m+wtSQySwhLE3G1T
lVNa9Ge+zMrKft4b22fPCcdGLaAJC0MmKwyAU9buzCne8l2fRf8yjHSAcpnX1L6zfWpFqEn4LsZ5
9MsIVSPNcwJbJ29gKQd5Fxqe7/GCPP5FQOxFPBbQd19wdEM5UkNe1ywUlhfv26U9GOK8HIP8o/xT
+JRD1FxhEfKTjle4Rs5CMwmWR6HQxF9PeGcSrE7S1zyWp1xXQj9EOX2QYOGDLjmHeDmBJWx0R5Ib
XwOUAf2o0Sfvtpw68wEmHsBF4s+3Ku8yCye2YsAYLK9ajDaNbO7/BkpPj6MWiJYqx3IXkhLDlXVA
Pn/9uKumJwndqQn6r686WQ32yIc5XzW18zxLE6AeScYrT2KlwLphC1uoff4e9fdfQt05p5TjmBqG
1v7TG0o+WG1CRwFVjPC7nPgC906JWibNkdGmAqSAewyOBQmZ9Q2/NNadJozEJGEDqD86Vs5cPELK
Rr30vVCsevX920YWYv8Bt+69AZHxq1nQ0kluhOKqQkpz41EaalLTpii/5TbClvmbQtus3FP5NEUi
k1tde5yo732Qwlk68A4eWaORmZeYL325ZANYKUl19krEvz76jXlO3bb+EMJ0UaVcugnwOspB08ll
cE2uId8Kyr74gAmc5QM+WEBL+H7KfevLH8nXNgduEyhqkuUjyqrFpGxxeayjPe027EF7GJVfyoYB
2LAkCdTzS9y8Awj3qr8EmHZk4GGdoyhR9s+pCVnzG4afv+bosLTBk9UXsRshYvXuL5sPCphYIwC8
UB316Iewk8P7Kj1jdWUCIzXj0mniLUmYKrCsFVSdR7fsL0DmARVmqBHbjKRJACG88AQtJU+ej5D1
El60jGSpXN32+gVUzI+ca/nq9RWkoQTHYatNOC0tCsue1dbPPPGEkNYC+PRszRF8s7dLv3GzkicC
65oVYAB4AQWxHpbKC36Px94MdXNCaRQO3Icz9Y/YO5oAbp0wNEMcGze1JOtJRbDhuUQ7qo1pCnAU
ZO/6FiQ9VaOr85uSAPMYVlMyFeeH8r/IC9I3FPSD/7cKXxdDrqr5zofoLJ0BX4PDXp1oYMbTPrNU
r/eFaQHOQX/vbB1bUKAiXonZCj5nHTXtgVrNrF7O5wfCQ8jRe5SBpzhXBYAR5B6/towlK+yXr0N/
CUEocEWYYGP6VWbUBAQeYJ5I9IYmH9EOFU7XcG7+jplO1UKcQJzse81mzd+1JqR25uX1GCsPR4eR
Vko9X+L8FFrhtdCYt81RNKkS2vN6E/yhoxAX/luthq1T0ajPvOISVN75YOeANlAegotHhpYGn2Bj
zuJLYEpvOPeGo7/xEUd4vz/rU/OY3iIDyJl4Myj0PPvFwGS8ZQvEG6nkxmP8fCDEzQFVxBQaTz8D
tyZCPGkzaHLhg2cUXUqFmLuPjiopUyDJxiEx3SRVNjWlwsyuMH2jsRcwn5mNIdcLTUKO4Iep6jFe
GZuQkGSa+evJj9xbKU8jTq9wpGFD+Nzd/Gz55ypTLMm+rcqgyphO7Gbz/1jMe6w0L2C6fEeQowah
V/Vv+4ea7fg2NIbaaY5f2+cYVPsO1p2JGCWc6DtZ2xUPg2YlSusQYBo7Yff0ESKXkcHCpEOKzfjM
StbFaJ0Ls+X4ouzijI0ZJ0bcsfSBSgsqIO1jyiqwR7PncgtTe54P9pb5X6VCtq7lL2r+xiY2ATGm
jcl7oTFz5at6NGwU08IlV/dHa58GxtCEOM4IO8e50rqNfTFBVWrgqv2r9J2CHg3gfH5GC9t2WLUG
lPmjDH+jNJcTesalAHpiEg24dCoyKSEp6iUx0XsTDAGh3ZEfgPg4yVnJtuCm1H7l/dexsoF1NmGz
rkcf88rilLbMDDrGpZOgYCUZL8BxlaAMdkercy/gm3HeH/LCWKSg/qoAj2rfIyji24Ye8buufakb
9lIWgUGPqWQtzry8Rz2XdKDaMRse6OHTwD+aDK82qjTpLdeOT25zLR98zwh/C30XMVRbPfMJrPUq
hJZHlDpo/ZMvgo96LvAQRJgtTMojqepy9hVo1VCoJXlQNDCp8VQtj4Sy977htO7A4YH2a9aqDvRy
TCa26+h5bOuZSZ2kMG+l9l3hlr6IF2EYHHSzcU+At8S1kyecBL0Qw617AkboNEE+bStBK/39vhPF
C9P14Xb7zSUIWnd0z2fp0pc9fySkaxlnUtfW+9ak/pjXefQDA9YgdGB8PVhiEyK/lcVY/N9UhLci
3LZZkB6Gurr95/FVK4L0GcfV4ajOFzsuoMEEls/0txu729ByJUkmDFsv/ImqVCQa1YhMG6wxrj9x
hAiE7BIHrjqei1LEsfzvjuCKzKZS+Cow2ZuP2HLFEBUGYPwbWgtgBZ2Bsm034A4nWPZF4RSOBwhk
L6wEGF03Oi5Ibvntrjkxb5C6rn01d7wzdKu+xgyOsdRBptNDbMu242JC5kdspEnu8MaGwaYcYA3c
m85fv2pmsQHr4lg7wo1lawzR+JDaChnd9IFM7YifnlUfnWQ/p6ZR6nFARRZHUl+9Ns7r+12W5i+Q
rSmw/TOl/3h8SL2fIUiMkbHZcSXd61WxwQm8CmGVYTNxZ7Zp+0W4TCCnWuUZSEqsoJbFvmUkRE2V
xEw5aVCANiKrgLmK/Wss62AwUX1ul6hirAmXCo2gtjwwLEaM38WlKkNcQjL0+UKoYJ6b51aueJpI
a+3ZWFO/2btA6kGkxBNdAE6eG+C1J63equFuaGq2u1IrgduTg2Xldmx184E//54DvoGi7oJnyk+0
oC4Rbrh44tUHW2EhCfBnFtZT3uCFOLjdQvmWuHel4T7utEXxjC2bJgHRYWuFJtOvAzig5f+tMXwm
hUk1NzLLHjvHox4mXphIkrGxEdJK3Thk8XZ4gmdUgli7j+uINUPE8x1vWK1xNApiuKRRWYZM4t7h
JT4ZKFrX8LuhPVlXuusIsNgrUgCNnBEXJRdkGiKM6zVq+Qwpi4ixdcCIhkdigd1wxTUaynYsPPxK
B4qdG8s/rHhJKCjuewem5cfXvkuraefzMH0M+9NjXVMLBr5Nl1ALl4XzWA7+HwN/874sRTyvTpOo
g7wzHgg716XA5mDNxlM3RRoXpQc93G10lHnsuqnOp+1rOgN0wNiT3XqZaMSRSle6Up+8aCa5JtJv
pPLfyNbkTDetzpYiHEWue8YqZzv+LE5E1USFpMkclQE5pes2Lqooo5CCRuXHl93+BFu3qInLiri6
u0gFMcuEzY/IpBa3/uHy8D2+weD6iydObTD9caMC07/jv2SRiE11SoN6+ZbwCl+TnWXVXzjXN2cl
EuymcS7zfJWLWOQ0erZZ3eBGEpcYyRfTqnKey7E8BgKALM5li3B+VNZL4NXsr6r2C6OlIYi1I8TM
IanKXCYHJMtqf1vhG/3T1Y+fwsogDw==
`protect end_protected
