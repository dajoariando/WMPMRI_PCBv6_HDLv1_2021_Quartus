-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
S6S98Wloo8e8pZqhyQFa98/ypVkpr7On9IgDgOrNjEjTvKGbkLzWdG0twolXUmPGTfGk8DypvNRZ
ebL7HuWbcLYlpyhi0JN5M+ZdILn/2nYVbiKF45bPKlPfk/McVts/xfMCGjfYHGpapEpmMuiQH1U5
Or28ds3hKBp2QfgpH0CzF5yY7w4ly7VaJFeszDbwpU0MunZUEAptGFo7/5k6As8gpGz0gdq8AtSN
/VizZdiS8aYwY3wO5LH9wKQPZZLXqqAqilIqRbjWyyZ0hNXYMJDwUZLa3gqgj922WvNuLEwBLMOB
15F1yJlLmhEGd2TV/OQvUJMSJcOkjyPx4nCnUQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4288)
`protect data_block
cutOK0Xc6EGV+z9guwOw9SKKaPdcWY+o1C4e5OFp75eNw195+nqFrfoFZglU+EyJbC2T3l5YH66q
pAEsjXqoiV9J0zFV4Ft7Bed4UfN0Ni7wAYPErNCWhpHLhCgIRAK+DqHDuhRA5nvW8k678kGVLddQ
oBFyqS3Zr3XoMqo4xzDHCq9xmH0d7qE/rLqh7Vn2NmOvnKeIzkUSSgn5pmO27U8TAJX5bbD8WePL
Vxn+4YpdLrPIErbUhaPRY3r6DRE9vIQ+inpElA7AKxARTM3gTAe/wtPfkveJGbOp47856sCp7Khb
hsAjdJfzviSu3J47MpFq5ErtMM4pgPdEilsyABzn5oJPM3aKSprihqLBSZAuiCis+Q6S25M1CElb
qNaz2+2lFRhZIQmG0afpY1QouACg/0qIGES0GWATtUsy7r+LZqaojlv080Y7dK98nlmymeQYikP7
N2Cc8HOdlTyxa7ndnf6prYl+O2ISz+9ZnYpkeAjLJ/IdwAorCbl5mJpJKp/r9voOHGGN0Gn01C9o
ieaWigUTa064RJg35TqjgX9YmEc0z2VR3v7EFza+iSr0Ns1dAkR4LsQjwq+fP/q2O68BPLVFyC79
2PfBYWNeOL7QTs9Gap4RnEa2ScygydnkjvsM3PyzgOq3ZkfzsymFciflG4E+JKmevDcaobT9IyM0
8XO0u5cNin2SE3u7QoN0InGWIeHGCG0DkKQGUG86IBb1W4fKB8k0/Ci+qqHzjl83KFGezOTiDNpL
Fts0qN8zZW+gyEN+c8cbK6n/Q5B4WNxoQF2NL5zgX0+K1Rig+PNHoOxowuq7g3fUpki9lTagIpnA
dRbqVmszyMPbg0UZTbKXBJJz0yr/61Sw6ipr0qcfogImdA4r+PZay96OwEMRXobPvtmlSjNk/DgJ
d7L2K8cNVzPEnSpt1G6SkQoqjfruMwRsGOyikTVEo2n373xlZvyl9v5B0fTxtTYtVcYC1FLyl8ae
KvrqBHVu5CpHhK1/nkBusO/opzFJbdu/twqmKiQrjDEmjuPcIX48eBp8lUe+lEvrajirOZLC46vv
bggy+qVBEGkE4/w0vTvQJVJkoqCSrbjWqrdep51MU6lMsBLlNFEwRMfKgNUwXAV4SOv5szA84Th+
YVn071Bjq8ojPNdgChOlqsThEZAIFVrZxIdeMpW+6hsXRfDqpExrA4zrHZjHrLTJUhAo+Pz9Tty1
cQTZWFcugZuwC783qVfs2QZg+JvDWJgt6f/t9sOCFk5C5H3QLAU6mblxwicYLlmC1o36xLnJHmM5
0wIE3jmGJC9lO4z+Trw9BqPB6QRElcGjIWv+om6y6jWdcWC66jcIULnN5klGH4BZn4K1nbgh/HBs
Cd1Wx0Nwv2DAJVUqLLepS1Sl/8ot3UQmDz4PHqNMcRh6UKwpfrTZel0Dl2rUY2Pk+dayQvM0+U9Y
gLULPN3sbvdsIGdNH1smYjg5NjiNYH4ivV34bJ93K/dQ5t3knYZlJO+A/4tLnKDJAvsyMIEKjpJv
pyQ+MWfYjce0815HyHLCWkPqNOouD5ujBwRxUSeC+i14WnHK7O5ZvKrmeZHhmaDq2GOkQp5YX9ZL
zIm0vf8kfJCsNODM37JHVf7wuFKX7yPUZv4zc72gb+y7TgRGb2sXVlqXRJgOFT6zxIuzs+0H4j86
3gBE+p6sUxoFni22wmE/98JORf0P0izU3gvWaewGJ/4u7UD3qMOdv8ZUEY0FH79bwYtjE+Rj/bDU
++wrjx0cuH86dkUwjZ9Fe/MkfrBnX5FhcyGLaPKhJCLZdp/OrgtSPlL0cIdz/tq9UsciepjCLsbB
dxaJ6Q8vWBG+eGTvlmZCiy7lTooXaXqRhLpPh0rKecDSfGLPaJE7UYkXWIQ3oorj38HiIS1HAlR7
YYgHRvbTTf5yYlNJEV7XzRtV0StvEyvJfCLchtNyiEhQRfe+k4I6ObpO3mL1y6h6iYlMvkJ4gABv
hf2DU7V+BLwN5ykmrYl0PXzzdFIOSeoDNb3/LQPOaEFhPhcWp7RwXGl0ozuSKpkiAYWM+KpqRJs4
1oK3PCO+m15tWqR2DQ5pFG/9vPryyODGDYCHTdYWwoOowZDo6WvmdE3m8mnJ1HShBY+fPt85SR0k
PCBnIwVbqwylkrmkMUY1v+w/cqY8DCto+mFH2HGw5RXp/KMAlG8YU3cUCJGgVv6pXkDzPZW02rg9
Cx2C51wjOyw1iv6mSrWuRi9J0iGuIode3RH5Am+xd4e5mdA3lI6IaLVAiHUDMpkKwT72/2zxIbuq
HAhXrkGOmbKpgFYwvuiWHXOdKhZMETIXw7S0MFHobNgWS/nu9/oX4yLF7GJBJOpG+7HMXEX9e/s8
akqYURFSljAlJxaCwWBH6HIUG1oI6csdAEm8oq3qik9oBX6kp48sA6cVUlNyS2P85qvQ+vEh5IVF
Wx5hvM31qeCMFmbbP/XSV3p7SpGHbRAfLFbbB1II6Ztt/+rLXjteZc23eT5b1bWMtsHJ+fWrNw9m
LzR2jTJIqWg2ygONWau1cqwXWBMsp+wA1umIti5RpstCrCrMzUTAy/0g628OebgCH1qJvAF1r5Ou
h5JCOXE41++GMyUxf0lVvjabWfxPuDeEiJ9NHP79As0ssUIKgDZmb8TdOcpaN6yvjmHBiFhe5z2q
xzmvqeHyQc6iPRz+MWTLxC+Tb4d5U11sPlJdiFya6Kn1YyCX/7a9YiNYd0z2otBYlytcAbwiPhXJ
nzAC/oTR5YIVRaOm4Uw+D8Z7MeDJXt/cD/KgpeAzC+M19arm5lkM52Y4DV9omQ9e7laSOtHehcY7
5Z+2UDy+6A4Xnt4cobLogttFL+7IEyR1LSwQ+h9dnUG7cLAtDzamoFKNUspAc1rqdnBx/mR0fhs+
3EQtCuWIe9FeQjZjMgt3cr3U23jW4RE0rvsPKaIekq1HShpmF2Rz0moergJ7GNBViAoYw739qv+A
D9oal17MJoTUG2PLfIT0rYqyxfDams6EN1O1SzjosiDlNsJHT8R7zk5EgQJL4ogG1mriW3AV8cqv
xsZCDnEYAe0yrpFDu9KpQ58HB9ZJmM53T2LPPiq1QK541TbrtaZqw/bmKGhLgPRsQquzgzsvvnNa
faHZjFwGBDHhlXR23WPRQtciSWN6FZ/kHSg2AM0VMH9opPus+2GR7nlVLAHmFQPmzlRHp1rcyUj2
/GbUcS+Z5Yk/ZXe0eNj7cmshXdl5QaYkWwCUU1gST4ZSAFEj4yz3QXZ2T/TqURVl/bJJ2yvL3GRC
OL18bbcy1vsyP+sy4k75B/8hwbOYFXT8rGNmZqEeXqEcTUzmi8AkZlrRUyXDrEt2aJEck7+KbAwN
BM6RAZjIM8eaLsxtoubtVPmhYgZg2AYFWygbg088shQQLJDR3iraogXlEUz+oR/lMeSbtG2sTNRt
Ml8GOTUSxrFGcGV6q6JqkMsNYHktCM32/Dw80Az4ihHfXrqI3XE60novfLZWzEmgBjoXL3SrA8gF
f8dpRa6/pnsy3MMjPpcW7jRO9wimvEe+C1sGe0VT5tEd6rfGNuYNVa9zOLd2/fzckgWbETgaSvUI
YFihKO98fkejEUk1BD1LB/5IgUUSaaeSxv6HBFcqBmx/tH6Kt7/z1lEg+QVMdnHsYKnDlCePmYOx
xcKYjnXjXutadOdp8+0525KuLMmVWeWeg0fS83bFR2MqzSRf1mnVbqI96b0LvWdVjAUPNmbmNZWt
BbsleyhICDfmFq7IoCHQs8irk2p3yTG2FuDDnHhEZZu1ZeQAv176DGoUK4wxXauFWEeSJ+1ALhR2
9OelY/iFDS5HZocKgDM0NpaTGRUPyudhzicpykiAsHc+QO/UIdxPy7J7y7fpCFVSEo1j/YGWXC7i
aVwHuUesjoyT79a9bNeyY6DVcbmj85+d1SE6nmlVbjc9MO3fQXXtbm/tGipEDSAmmWEnfdJpfdbM
BeBlvSyDS8cpTtQxgQbbzD7TlyDZpLU1LAAldkdu5EJjHnW/BSTg3AW8EsgEDYomHviW1cDRtMC6
p+vtlSnQk28aEe11N+MecEnBdaIUvix+i2aTXNZvd137Zvy4JJJgPY5dNdSFXVCRqvQ9V69AUolr
WsbzAuttDUB2LfeKEBExD52E1+21f/iW/mHyNteENFXF2iOh3wbHKSrRU2+h17AahxJGQHUCQVXm
sRxlM7tavZeSHmj9Etat4t4jzBTRtBkWruiheu6APkYEUxC69qwQ+ZShViNFOcn61eh65E4bMjNo
7xf5n2rqzyn9/uVOlQs2zANIwbHhHXUHu+JpMhZScSTA8wuQWjLyLZLrT8awiEG6PWI+scLuyTm/
yo1P2cGE0acuUg6d4QMCAMbUKklWvexcDCyC8LA+syXXpoYVrfT5fGQJFW89iOEr3Lw5MLqBfTxu
rDnGKVlWwYJ6N/FSsMc396y0tPFTs2ffBJsuNcnV5FmdeA56rV3nrFTreF0TTgcQd22oiCZ2iGtf
Y/isQw+vNsKNWTCe7n7bQbr24cSY/owqIwHikydzF5qhjGKB4pIxg6A+aYVPxF6E/pBCz9KwsosI
4djDWZxQNoCC+WY/eB1sh1c7IzobgCFH5OAmCPcFA6YzVLs0YWTTSamDgiZt66cFOM2BILntQkIu
dSU1jT5ZcpRzamKiE0uAp7EQYbWHkCzzsGzQhb81qf4rWaiW4LvE1j9PZn2hDWrm19hTsLJ5J9YD
rQtbv7aDc1rT/tqGH4jAg5APWvnJxyL1JPtfvMSBDfKrv8gMewEgVfdF7AWaW4r3f+B7qwstvnKP
KpUScf0SJ98foC0QxWsgRPVg4OuK9Lggle4YWP93YnxGKZBktgzFhJF9cXm4mm8W7EKRhAsFxIyl
q9wCbJPuXgyvZoWXTcfjWqY2sqnHJOr9jsF+scPXWLhSQ1TBOQHUCKNs/cPlwfcWopV2uAw1bCHQ
H+nNzEu4HTgJDhCPYOE2V6mSaSgWmtifsfPK9GuEtFFRzykjiiDHyEe09uqwuzCMzvWj7VpFnZEa
2VEhcZW9UyhZhFKP6DccA25eM0YtaNUtdWqmh2plbR0F50wUUZSjg/1eGgW3O9fsXkrcKf8d7qf9
B0Y1rJon3XxMuxRRpSRDM9HcaCMQuZNYNGd+MFbDVROvTDnwh7L2KlknX3ovVIvivwyFErkYtcd4
uyADHOgukoyrfqfD1h9gu3AKyV7UEwUmexYulRz6t9zPW746OKhnNv4BYdsB7eKarH6DCyHeVZTr
zo8wAdHvH9dJpK8qYxjzs08uK2yA8u1qSOG3wGX0HcH36wuqzMA5I/vk16oxdyx/VCuhdV+gdhvc
/P9VHMWAif6qfilZXm0ach1DiusB6D4XmnWA8ay49cCOPPd6kI/QD79gYTH7Twyz9URnIztfftPa
XCwTIFBPjevkvIoYovmh5bx9zPdOp1NTysHgsAm5t5+M/v9g5yJGLjX7G9+VjrEq3f94mOJ5m2cw
CB8BbcFi/ZhQeJTjMGRhTEuoNK67ftyrpwc7XvDU3kKKMKShs+GbG/C4nWGOo7Jh4hJ6Ll4uUfNx
c7lzi0kPEqkyDWRPsy4rRr/+De/Qtr2/svzH1vRkps9tTS4e7042gcRYayZu0cR1dgBPEOgaj+Gn
aRxO5yKN3qvbmT/nGiwo5+4gi7fn0E7uggHBRXeo7aGt9KczYAazOIRbVApwvzo5mu2yuk2L6nVg
gKrwCrYO8CrOvJdP6A==
`protect end_protected
