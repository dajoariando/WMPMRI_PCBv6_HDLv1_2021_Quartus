-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
AY3QKU7kdI6eht15KPgC8JFi00kpxBLHN+0zwETw4wqj3bit9/1KFt3Laxgqs73u09gHs30nl/Lf
Cur+177B+XA5DDYeo4yYAdZcLRc5zcREtvBcescEFCfpSGBLgSBD5CyhaAlDzp5LoDgBXQz6mrLx
LCbgiTX0d4yTIAu6sq8MX0+oSxh1A/S+4ar9tRVpgpQSD7lEXQCnzvzUls6XAwF9Kx0+nDl9Tx37
rXZAynZFSPVT5eG7RlNVuTOzNhomFoDvCu5DqbQIx/4i24S0ucamwfLOvwFYTKckeWRuFt1f0pbO
bAHI4Kz99N5UOJDjlYoTTCoz0nYCcis7Jdu6Sg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3024)
`protect data_block
7tbfzKokayYaFDfu7VDVEbd2Zh10SPYN/RfZO2+7IOTnba4j19/AKEOpVjtKYiCMkjOirddO2vki
/PFpr2rfKf37iWpy/hmGWzBCkSx3bdTwMY7pxNtfkeu87tpZ6axNt/IaJyrjuDfF1qLMWIGAeTGg
oNYFUzW/eQaKNzun6DQPq23N/ae9NO2szUOYpb94HJoWOahE1H5iYbxpwg2Az3ZF/3ihFVQcQiPC
vINUKTVEaUvdlihXHl1Mt1MV4qY0MqZmfD3Ji2dZpzfJDiwgbtdwqFyunxjscWkdFMXBDeXBLgdM
drziWw3xtsRhjJFN6B1rLF9x3hwJD/BqL/jx2V8AV1bL+u8zbHY3+EXXi60O64NRHB0nZxxtG9vi
saH3+xmVHhxTpPu+WIXZOL8YO2tM/NPckFUvj9tCnTQcniGtSVmXRiusdDYKScXbLF2FBNkZsXRg
6yU7EcEKkqTMIjuWUO0Y2xKgqTdPj4uFLYG5X7OuMTekstLdhfMNR6XGLnv+aPtneuyLAxl4p/9i
Fth5rPJATaFDA6ce+4JZdbt3JVkP9/j6iroZcv9r9YRC8b0nWxnDbkB8+XVt0R450gyANApqisvo
Hes3Ge+TQbnu7D75A2HxmWi88vBuIecNkf6DjeaaPx2BC6TMnifzooKJbtnvnx4NsfUPsz7aJZkA
HW/4O5h0apt+EKoIIb8UJ9bY0EUdBbbTStd8fCoq2sCCPvc81SuXiRQcfhOPvwTB8Ih7k8CIiAXn
98QAt6o0rBrRrCH1VxPUPPmuwyfI0+ceWQ5Lkq10sW5S9i9OAVwbsxZNwVbHlJXf7kGy3lW9vDDC
k4kVi6sN4bAovDIYXkEzEQKU4NfSfBNqgl10xmvbJhQKt+K8oXT97K81AYvSqp8RsD3zbh1IU5VS
W9SVah0XaEZwRCNbgNSg+3KZtm4n8k6/HkGgUxmIiqupPR1SmR6soQlSiDhlK+/HcnwrZPI2hv8B
1arFUH9tCoeTcwqyWI7h8Qq6JtOKqOdRcF01JLhrgQPBQfvb1ytj04eSD734hJwuuABW7agE1rLV
teb/Z7UrI9vhpapJXD2zNVMhwaf0rMpKT27JCyidWuAkacKaz1WLRASQtMuZmWZsrncnx2V636wM
W7buSQD3luL88joozWGHNiehjlDDZFFX4WwhGIyNWO961uKuH2PAf6IIfvIwgmDFwMsXB0BFi2x8
HIeE/xzKtsu+ycgCO9GWCpkJQ8Gi/EcqarREjMv725ONOBbcnUnNv+QA1kSG8r0Bvzj0juaJggba
rDPtGW8NAy8aAyiKWrAIG9eDaEaS+fKTsLYE0NLyrdZ5EJO/s5prPDppK1Fljnw7DasV8txGS86M
ZpNFGan2463DIFys3Gl1+hTLvK0kxwzBIAZEsA75kvZXXVkn9BU/DWgUz2OQBoFIGCywR6lgiYZv
b9Z1iGG42Ov1UuCpbzK9++50LOtxUeJfQN9sb5q5QRcLT9CBzFV38HEP5mWH5q4TbSjC/HnMXCzf
qpDbhWZXZCUn2Ep0V3GCAc8gA4Mh7rm5ilCVbZ9Lp/UkdFxXUYHL7IoLgKyizsEjElHpreJIIg1D
cbH/oH6OhKh9T3OPMd7fwCNDNqm3UE6sYqLvQe5dMH0qI8JJvcqv98cip/gMSNSfPZgkcnvf23Cm
BPOl2xfStQn/qqKSAkPPgAb5EmuKHeh8blbuxeTmXZ0wBxBlW3eEXRWzY1cWcoJ779/0954xCWi8
FnjAn7FLHDMroD1+H4kGfINQZwVujL1U9V2hz+aIaOzX37ibjVx4DhSrsy+o2wnCSozmbdWenBXT
2JT7w7OwiEdP7vYtEQfsiiEk84UrQZYrmXWG60IPO9aTfnzdWxN8BisoNrUczL8GPz8EoH4wQMfj
k8RIG5WEIuea7hKUczmiG9f4EL0tu8cHEVr/lb0vhIX8hSDB2UhtNMcGqezIJS4PsEeoVbJNa70Z
Fpumo5HY2rZj05Vi8Mp60zqeF6kzCRwb0yOBnSfw+C50Idz/tDehF/z5RmPIh/Ys/rNiks4qV9sE
i5PCTJu3GRRWCIWp75oaV6E9FPVg5t/fs7q4yYLR4dgeBCi92zf7c6Bc9BrjDD6KvRjuPXxdR//W
jzQhYUSGCY5H55VUxE4NheYBJyY21ufnlx/O0yLX328Bnc28OC9NTg1/lp0t/A0zvPk37h5ShzT2
yPlmn2cnMSsPElTDnBGUkQourOb5pSlgQBoibF+/PQ1s/ObLTs0TY76FFwjAvRua+K9qngJjGDYi
TpEOiTgxf3qzHobqepOCxK9+fC0X7BNt1aKymts1hGMR7fBLHUJ0xfAVgWRzALndNDUnMkOaqQeX
n9T4hr1wY1T2/eqOiJkJ4+4kObjgHssHXWSsKVpxdYsjkFTzMgudnwH3B+Lo/t+x7Ypqb2/sPt/p
Lc9tX2B3VZ+7PbUwAzVc848Q9uYr7muZlUCvUHtUXTZoHbygIbeZb9qhCi0zFg1lSJYzPMcCkTFL
jAyoQxbOI37DR59wirtY+RW06x2JHF9f9UPWwxHfYIw3QOxOY/na3k8KSB0Y4bEoSbFhDbYruCRw
Y9ARIhJ1ygJIeEFvAf7qhOe/0ypbbhdP6iFOH4XzzSOw9ziQyuQKhB4SI5wM/4pS5toPU0z+ZaJt
5PMxnO7e6yzRjqjjNq6awgUq0vbl3244Yr+0fZsBC+S/TnoMUchdie2FXsQZF/MEtNJtvk9mGj8z
VwUNCsfWNn6+xT5QRtbhAUxJdo+pALXtK7Zhgk2Q3m4rTbU57hrnM9ozIIuSLbjnkedUZRZ0cn01
dgPOJ44PEk7ebsoMeZ7QlHEPEai8h+T5KPDrK28uT0hAJ2CCtJbecAxbRvWun6bWeKStKXpTUWEd
OsCMrybK5MbprfhS2RDYEorM8VNFGY4iPcdw7zbapSed3zLrLN4H8IrEaZymMEwbOcEWDOo8A6fe
ZuTfP8Pg/HdDSh5iSUUnsVsTwn99M8JPtzvPGjBC+nAoaRPSD5u/AOkvSoqwN/VQbMOdPaEZZ3X0
JTf14TuLCwGI7Ut2AWWCSZ7o+HdfemmpWuBH20XytdMtY4jUtXcB4UCo3UXsgpyvo7vHMA0CjA00
QdJesrOESFPXBICUM6EFv0lBHrqyJVorauWQGwENN3LFnK6KtehOFtH0aImxFGjoEuNIbneBjKB9
jYL7gZ27o6ynAzcK2JyW58pG2Qoa/IRXpp4loyRObsLS8vCmLCIYgUMiSJAONXTTBubJscRHOJte
ngWiNMOuJ/3HGQeiafNS9S4ch3K3CZAqlQIRFrsiYXHGzJLjJ2P4eUd79pfvmMn1H6fiBi0q9vZb
fbubnBnV1T9/mprNyQKwa5rIhITH49EAcqWeACYLo61hKAAdpoFmClTku0fflnQP+ERj8d4Quk++
Eo5z8zlSeD/Z4J+1Nx7PvWm+EdDuoatMvGxbTKjlivpsXUelhydvXNvDPpI91HihHVLnLOM8tEVk
ULUwNDcKWqr5JL/G8BSh0EdOOsDj9Ki5RG5+vYboF1nXy6K6docg2uLbmdWCpmFAC+9Q0y5P7UR6
AqkE3f/oJnK7Dop2NPLlm0yMEZse3qI138sq1YO1fECm6Dhg/eULcMTXEFYnqupx1AeOx/jLWFj/
xB6V6L05YZmsJtZa/yNjtuEM1KLksNGAa5ZcoX+Fh90M4724yrpxyPdzGy3RACXjFZfEehnRiNg/
sFv9sUO5nMtHgmbTaHeRWQiwdjMXK3zhye/FZOZLmnNwxExL4HrTNLVRlvheY3/rlyY5MDW7eH5w
bSFaEf296GMqaLQ/UhGrEhTniVyjHVHxz/6TZft6YkUS0o/DsIY371+rDs1rfiRoQiO91gmqXPMI
TbnEBob/xW0MxUgziiwyFzRC6RDnbcEOHGBERGL5WcUZWCZZgsz+BRrbuIBpX/oOqPYPtqubGaJT
lrvRoxx5U2Cw44bHVbsIVPhQ4dd33SZjH7kFJuZQ3It7pRgHz583Bk3JEC4rS5HCcTkI++HFNzpa
cJdA
`protect end_protected
