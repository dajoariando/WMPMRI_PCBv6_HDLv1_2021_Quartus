-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
eT4k7ADJwTi6qSSFyEdC4ZqGESEcXdtZVzUmb97fnwXdkxGGrtlLeqhlGicxrGoaMjvDd0hPS/hb
LyLjHAS/hsYAIORzhsWJ4aVyqhM7G/4ACL87df/t4mAvcDSGyIfHLcIrIAuKR0mzmVE08P1GFEhQ
H4fN4vvV9N30PPxWE14JGRkJKhPzXia0/Mr1dpyUoFQD6Wh0S5djIcsZzhrnIyRlhDvHoDIbBD8h
gInBWR199FmbRtZS+vioBXXMt9c2BnFyxgjoJKURyrIu4SjWib3u9h9b1UI3+mXiY6pNxlGmLTZX
39A0ThZQ69yjJAY1vSFj3G4bvtIinTijhtzH9w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12384)
`protect data_block
7aL/Vik9mbzlfdyH6floOccW76+7DeKcaHPf8ZwoTUc364s+jCcLRhm1x9onjgoXxI1o95DgXkUi
RzGrI8UxcqFeEDlPvdERqhNplW/Vl1YFGdOAgqJlRg1SZzoDGUzcRvqnJmvH3prBMQTo3FZwkh8n
l3iZRk0E8xGs3z79zwVpJr6zw29U3GDX+DO05GysWptRMr7FLp+N+8Icpz8jwFXsOv9cwyLLvHM8
+3w5a2hQJq/6N+w5WBrU3qj0LQxvRIaKUmbdnZ1Jun2R95ijA+4VKlqJ45jiKd7Fv3jG9zCYHnyn
vttJ6YH1CvkSi3iuUY6s3V5S2mhPIVCXMy9ZLZHgBTkYaueJZP7MIDVsL9NMZsr7sDe0ygBGmaVs
L4Soa/UAZ0IJ4PhNLAhtF+oya93PxcflK/sBpBJe0mtIxYv2ToVvB/FVhrQrS/vaRM70R71xKCeW
cCNL2eNoayK6DOAU7RyW7c1+lkPBGbJyRKh3D6ohlQ+lDm9+VXs23jj2p8wevItNBUFUntffn0NF
UHnvEGAKIjjNO5LxnQAc9n9RxUn/iyVrd9xSV6T84stYg+uk8CkoipoUZsVhEBUjjV7No3un7LOd
U+P4VJ5nr32BaoPXemYVKJPZJAbhfP5ZbFBTF7oJIqxaQBUlo847DfXYrzLGUlwcoTQNQWKc9DF0
cqlqauLweEpvRYGHk8I0Johi1fBH6JpXAa+kTyh4MEAB5hL3ujgj042UPpHLlDybrPcQZbzhA2Bj
tuHEYTr2ZRwGGoow11XmQyczckmafYJJj5WCuFEKAvpcpfyqhzQ64DOznP+pJp/doeVU+d/bWfS+
tz2M6Cu2gmfDm0wgO/7V4q8vMQhLNUtNGGT01/RT0pK8ASD7jaaUAhDBBhFxTmHx2E7u/udVOSHD
E3Akdk6YKWvqXe50BZmPXvPFSZtom0GBUCi4uwZJedI6w+M1Q2nYrxFfGBhkLYNu/3VXoEweNubZ
hf/6jDhmlgny9RhnF8brw8br4Q61o80srSIlQAm2cVNqeHw/+StHoG/m8tggg9u15XlFNfZPKwfY
bFHeTpZF9TUnBoChYIu3b4copbYuNlrLcgvvQ9z2h3ChVyc+0EiY99qlvH/H3sLeNpvhkqw6y9d2
E7qIvatmy8o8A6OADUiAI98vzzdoATDQ94/DpF/t3cX/Bs2ImXFk/uXt48HbdjQeV9H4FsEtMiQA
57/y2YSJjR8jlc1vWof0XKYQytvslb95cOrIFe225iqJsh3cgrXeS+fkwcW0qtA40hKMBl8Y3xdZ
kCSfdyYwD34iYx5zDxRJdh9YEAVa4c6IOjTKtB+aF+cJn6WljfLHTRmlLUJaqaiQYdmiHE9AStuI
zx2up8+oeayIgRMPMsdgKbN5rwlL0LrCx7aDXpTWKsIA8bJraBd4kwpvNh30GLRNepBWnK8o68qX
DwiZMdQ8s9JLbzp8zpv5wtVEJeKn1rxvY6aS69gzyvg0oAjjp6GMIt3+OTulg7J9fBjJbR4lOh64
216lSlBwYcidb1IJ5ic+d9xmDhrmwAYSUovdlpSQVy6gpPDLygWRgqf/uILsYZxxi/hSA4l1hbxt
16Jfc8hjDjWb+CfANz6DkWof3oNGdEAXqCmQqOyuCK/Cj8XFrED/iB6ZglJ0qKtfKjrvseauZ/YC
YeZMtFUmupl0MuxOvPy1Vck0UqEyt6+kahKaDVKrzrTb2JX5swbjVxEZjiVDAKGg/0QH0u87UEVW
slhG9z4EdSxaNIpYKeJ2Pi9i7U2b3RMFQwMQ1IC2dkO+XmALHQihdkO/Jto1iwYIXpcUNJPiLYhM
MRAKP6cEr44LAntWdgbVbxaBvlSp5+QPU4VeVJizhM3FMYLVae8OripyFMqVOeYfO/fcDA4fdua+
ATocitozPPt6R5p8kfmvmgivAdvWkeuZlI41lrugaycT1Dzb1gOuO7LKghnwqFHfEVO9xC4PKaAy
UQzP56GomDZKmEdtrtoFgz34e4KbZIoC1712njnDTAEb0aWbN0wugBs55CWPJGhHiQ87vgtzfaOh
GGJ30PJYBI/jDXFSTU1XWfEbjyDzFC1fTQVyXl5pALD1xwU6aJXCTAkdDfWCXVf5QYjlMmcWaGkB
ccw11SfbjEC4zGcb90ScDXBvJNvUGiyKMsFz1KMiGL5jDfDT4fdH0oSmTYlSpPYOw85saUEZoE51
dLX+OSoz2/G2YXa+UxWD23MXtK4ohebwks3VYrgYmBdsIVoFW4Vjyfe+OKlPAfgxcX7nGoO6kz3H
0xc3zvQcDS5FU9x0QJppUzPuzN8FOR0IBMGH8fZycbztBmLz/+jVwRc6YDziaBpweJBgLyFMrcDa
ag9Y7jX4AaTZVUFzdEg9cAt+59TmNAHZUS6OhLduxhPsPQrXj8g7Y9z5vChgrYIGBNrFCHcJ+Ulc
k3dl/SHUiAVsgxEhZ04G6Tsm95/UtKvFS+iEXUt1aztskjMAqaRmcokqnkg4HAADJWx8jcgkZYoj
4P2VJLR4TBoe4MRrgiAgVartsiJ/wHRhc1c3uBTsg92ZBnEz7C7oKc1bBaozrhoMaztTl8YEA8y5
KNSTBTQ831QaIQ6DnrTKCxyzfU1NkqXKv+BHotxgnun4ADzme7tAJy4Jykn3APOp+zCR+jaWXKVQ
1gDlJEWjWAktGSCQw7rQgmnATazsLcu0ZO6wIBIZrVlTtHX5VgRW1FZYUCRua+TaSJgEXUktVFdG
t4FlFcP69BVUZLej9FS3yp95xk5vJq6C932ci/5VRwwKadH32UngloFuzBt1cbAJxNEpShfnBEbd
UHm2tZTlr4AqIFu2BTEUUze38gSr0K9zoNNEIHp5YJl5Fc0vu76m7TQEApGQ672AOWuAW+PcgAc2
2UWjSV5/LB+wm/Pio/ogIMqYSfaiV9ZM2UXdsOJkaLz7oKMNRufN8DPkb4K+B/Plnn7pQl4TqEK9
Jn1j8Xr+SwC5mtGveatoTFflipSYp2fZjlyQFHQ/XGSAsaKrkf6zRBjqjzcL/GW90eD+K7veZtEx
EWZ6XYaHEnG0F93n47ADpKA8RBYcW0H7W5hNME6wxw8UKpbZ9qFM20yDDo1UFC8IEnGcFD3+4Qjm
3wWPHI6XIuI6Sud8OHkS9l0z4lAaaiW8gjs3oVnbP4myWPfu1O21MDzGwoHnihNY5jE1KWldupxL
pSVGpVKtVn/D2x8OgtPK3X6oTGKI2aQ1hyicb7CLDZiP1D/wsjbABaM/armTmuf470QFnCcxE9UO
vnXjFPwAGrb3X+iyGsuy5lwWiHH2JDbab31OqeBcaT6+ke+8a/l9h0FvWiBHva5G3K/iYHEN2UBA
onqr7MBVDola5iQBCMMmZEx3BHOSL7VUZW3mPFoOmbdxuNI/2PuuTeHB0YUcCKb8Hbrsk+Sf79Kn
ADdF3+9c7pNZhWc2po8w5L9Mv/wk2K6dAd7pW+BRC1fgatStl/Th9BXaWNLDfdmf4quofEKh6KNo
TtD6ysnyNZgNFllbCC7ROy/EtK2owxlJQH1u/8y3bvB92r2O8xAluYTZhsMWd6iwW2H8sAlUvgaX
Cu5hNgV6/sEBriQ5E+qxtvwgSU4WZUqCX3THLuYBRX0VVMYXKbn1vXk3eRh29aufXem1mE4HXjle
DaexoUkbXH3i/jUFbCQXif6p0Ln1W/SxrAwueai8bj5OLTS4FCC3+iHThaRwPyGHCAKRhxFLPR30
WQ/7bFf2Tf5VLpoXyCevtKBuW8JUPwl/CPwHUJWAtgPo0MnqHBSWVE5sMTYom9xKgPgcs6itPHgx
T/2q0TA7aJnODig9XXp7aJBXros65Mx1kVTlScAXJJDofzYLHov6hMqnKJGVwM7TxwVS7jMS0CvI
8zkdbCFSQyDDkf0PKRL3JHUNlnJgiPVh7fMRsH8AaBzPCJxY6QqxGSyF4qBfJYlNYC6LAiWRP0u8
MPsMoPgdjw4DtQz4xc6kcVCDDPkn8fuPwZxhnkrlmBxZe4VQos5ytHshaQ/JFYEJQWgRXNEvzecz
mMSGTjp9giHFVCpR66lqUOB6EqlthSsC1GO4JdAKedI7o69QPjG4u6MJVSM1Uwg5fDvY/t/QMFNj
UW0X54OG8H8g8lvr64k03jIr7J8whoR81qDxJDDBuCKvC7v1mL0TdHqyY1ZtLY2vU2MgSfl+riwQ
nV7SzwgljrUppQ6cLrDaFHtmgfSF6z5VXveRRUBcD1CV5G+23CjPCz9CQtOM1WzaV7KusAZlRdyx
Lmvpm4ZZ/t7YgiMxN9vgOgRPQ/tc6tZehpcrYIMLOz0Q/3Yu13bO7M5lg5y1sAL6aaha2J01Q7Ud
XZcj1FMhk9asDvCcO2vmQjDQPEpJzV3fL4jDcVQD5ZTL68Pvt8olEEz+S65b7GOBFgXNnS8IljdC
On2BMyl1nJl8m/qWZ9cbEsQsNn5HMm8y6PXQLy7mZtGsCIL7qOiFZJkdg57NjmetZ7fBas8k+dvc
QvWboTVh52MU2lIRsMvTVbPTYlh6cikk/JUZCBifQMJ460wYxl/ey4c+K6iPESdJmvAkKcohzGBT
8t+O6YDnia2rKhfqHfIJvZL4IHexuCl1k7uoyskduTrCIQLdGwqvNqNo8YQNqGhUfemXQhfjO2+J
hSwQTQZjAvhWIkxw6BsK8HpFZWsxpBjauyvDb5/rZ3csOrsTvShd60n/Q/2kvwgAPBszKUxve0F3
Mq8lhQ5GhWSNz3aOZhUt2Ui7OEcHtQJD04cvM998RAi9niChnoYbvpsFjN+UZ/kXmwPRSYfLfNqK
GFhKZn7wBSOZNMyhFnDrMe5S46gEeDNi+Z8/1NldON/MpBspBePJ4y8w0+vfSUyJvpIwjeuTE1nt
agYTeQpP6hw5Z2gp1cDDVy/1UJVbrSvLo6PEqUordB2IoYSw/r1Rg6TKaJ85AqDjWlSt+Q68FLvF
ZodMU6JKdnOsJPqWomconWCQ8UluugpmhGngFwsiq+AZnfxqy8VaAhGJaRCcH7Pa+c5lLfPUrJoQ
hvZIrmpy8re5YQhY8tOwo9jkS3dk3OdeNUk0ho3TDsopPy0lM9R8t3PKRfFUmKeyMglEFV6FZUd4
9ueaGQvP5WBGgdo1uaHi+ooNTgBrw0ILwy0DtHLxW7Y/Zdi+iBcyPOj9k3oD3cSnd0CgNF2yCdOQ
XedPnVIEWqENOuNLZMksbU9OoN5g//bmXuMsNa/sn9+pMduyWLtUL2PA4aSgd7t6VJrx+GxPMsJy
cbWptzw42/do2bZ2n5OlYeR9vTjxXduXrHI+V3ahNHC/KzcYrQc2LTkWs7pWTQbo3XsU62fh7c2D
pHRNO4b3kR2/T+riYwG957ZZTQLTFn397FRxUknJGMlcJUHaf7RhIQOUfhjdQyxWtmkIBkpt1nIJ
VR1a+3QYH/DgwQpcPI3BRZk9PnyXMt7sVZjxmifauFX+UbqK9zQFF+Toa9EK+dzVKA5m6AgzTXyX
zkT3J4axADZhL/cgx4FWsEXVn9WehWHun3T20ULvz5KTZBaIa/ggDp8WhwIPaps7xsPGLVpMX5Eo
pzeawg5B+kXAbDbPmk8FIWHzj1pXiQNXXnNoIiA8pIoALHUIwEkoV2jBNTyUSLmuCP7ZW+sJctKu
CjrVi8B8lqnqG5KAVCnGa4pobE/kPawvm1Io1d27gmrQTIovAl79Y7wSfMbS2W5ri8E+e9KLRp4X
vPvpJY3YILvn0j6TY+6kIOLcSPT78vDFEF60h/ai50jws2CWLaNmyvXnfd5yf26gz5bzKsCwYNQF
zyvyhAreFV3y4pnj/IkbjsKYSsfkNIR3DQWbMM1l8MHkrSfT+QAWd2UNf/uw3TblGYVPdO1Zqyyl
jy59YxwJPW/96mKXEitAvixxOK3bX2zZFuMZpMYaRVDW8bHPt2+RbBIB37uhIDTpKfUFyMiYLrf2
tx4I0jHs8kcKSxtceRgtU8hUvVQf6Wade6ZA4OhMmRs+OCJGpup7FqQgP9rGK4/xbRTDfcfsJh2G
eHx0f0W64EZEGy2Rir+7zcjxc7OsEvm5Iscq7YZnynDGiLrEz+TYi5P7vyA9BVHOgG48ZwaoymAQ
/g+xakMHxmhJzBXnFx07Qwiw3mf+mgNULQLS6oZdeM/lEY9foPYiTI5n3V6Qivr7cq0iwMuy4/Zy
lFf80URCNhtdloiYurrkgzfMoAWSJzJztih1p9ywZNlM9Uj/Emhvf+zqVB2Fh7KfhC+F4zxAwxDo
A4WrLlckLYcSQUmXsHIwUBSlMlf88bu7iHoDIwTH33wt36c0evr2IYCKM/yf7fhSUJyJ8B+eK6po
iJ3pn4HsghGru1+uHJTSaKnHd4YESFcgWVWu8MnfCttODHo836P/wkNcewY+4LSXfzC+sZdhsVqU
8MMsU4w+5X72qsvapwwC50TuWGf5KN/Xb/Qr7A1UICZt+8UBFQB+t098V1pd8AuqX2aWhHrNv7nC
xRtEuxJceCxfd/m/3DQ8sXSIA9wQjx/lQMIKrDamTbcANf2uBFm1vMz1qwQaiYq+48lu8sl/NcbC
hDGgj9rzKqkSrKwVlPkZl6N+OGXSWLS2JZm4ioTCNcpr4iInMo7DlvpxypeUDxMPXOHkppf+yOdC
ahyGeCYpwFE80bfPt2tkeON3OM7u7zdE4tGrWN5uHdVxCN1RgdZvXIgNMsBMES4/2b0qJNPrWtJr
WvobUuyWCu3EC58DhhE9HlexWhcywYJbaZKA3wxgR2knp8Pg5U9RKp0gEXraBqlxj8ZzQ9Sx4xG1
qDWMXKmc2hK3EbpR3byRlNsg6IxKDEB/wsBLVRnGEqmMBTcXA6NrDRbefdrP+Xu54thKcuJmfQxV
xzDQfYZYizjcKbOhZ35bX6qMoWLV6kEaA8xB7axzAVzj6TZtAbX9rVKcPh12+x8JahA5XNUfbWG2
Tm9k7M517qUlHOn60YEXyAxzsE6c+IT+HKfap1KtgJMPVrNNqI3Qm44zCo14X7jshSb84a444icC
HsGCvWq/AGnqgRUAcEAWwXC68Tq6vMIFBJ634voyacegdd+a6JcTzQvl/qieTb5RZDx9HnPlVmUm
vI5MXGcPeUcUJe9ICTnt5PgLJwF0H38O4m3ln8AdlD6f6kU3zz1ET3UqbGbK4pUX2fXz7HaztEO8
+3579u3gj3EghMq+77GfAlJaLo9ulT9h7pI7vs5T36ZozlzMfckQx0lBxwnKlmkNp0QYhyepUD+W
XrXzi/2eFbY/vzA+KOgwU+hyOYExYveCzYJ/ViD4HRIw38hlB7HSZSyv7BDdl+x5DveDHgALzPi6
bK2QL3DFbGnfqdMkIUxceZKF9ZYi1Rl63JZEnZZ5VZmcR/6fxtJi5ijzQN2EYvV3fV5bOe0zVHSs
LRE+uRlTIj6F+XZbwK2N/rynu+41ywjev8Dsvas39u6SSviaVcVVO9gMu2oPfHqetdrV7fekLkTu
aAAPiwlq91bRUgaYVWlgk15/pUi0DHqwE6LcQBqvXEkXh0oVNrlWlg2whB0I3Gj2d4fSMEBiFNm9
Cbn2c6BhDOY4KuFn/XV7vcUb0bBWI/Xy1MwqeZf3g76/QoX8dOJTPNISVzJ/l2oBzqvGAY72kOav
/iW0MtZuSf+kg0WZQbPG+xs1UJHc5sPzSwGRD9y2PlnsLj7eh3IWnfMKdOyCknh52BxRF8AZVsSr
9WtFyzv3yZ6415F8ky03yM226v767ZYIVFKBcizyH5Ku1IplASSlzKxPsb6LvvI8juuDEO8wAAa3
cDKnmBJf0CfrOHIjzRjQsz0we/zR7SJnxxsnVVCIKFyESoOAXUvg4IV98LvZZM/T8wXTWTeLGi5J
2PsrqWitAfk3feqBcMnskpDCp2psoyfkPCFq0SDzJMsnvNWHF9EJEr9X0N5KGob5UxKPNGUdyyTc
4VmvL3Q8Q4HgTkOWGHIb3ishie/3bC3bj5v81DvUwH4x/6qWMnG6kQdSFlrvYGHkkhQYg3ti2okW
HZod7s5aK881Lh+gUmCL+vs6z5+9MhnEjK0ZheF1oqCz5Z/240E4bsCtNtc6gbIkHOUmdu/3RCbh
j7Y0oVXwlBD5yFbFCalS4N9hRanIuo7R4Oir9UtHKT9VpWdTCh79eJfnPMhlBnKUucXHZyyJnkOc
0QvAZMudHV6+/N7asj6RdQrg/LnnaFBJ0ZWXNpJtOh0yFbkr/vRLxt6FbfcfLzSnZmWxS2UTh9so
IVXCi8hhtbgVLA3vyXQBGK+OBTCOjefLjA7sqA2Sh2k+0xDajzRRA+6t3Qh1NXlsxwf47V8bT4st
nwSCPXEWTCtOqqpfIy3w45NAQDCoRzKOBy0bkV4a3AaDSngaUIbGrsR4hHLndq/7ZYdOgoBkIDcy
ukNSYNMBsZNwZ6ZUIII7rSbtiFG3P4h3bS+UeIlFwaeLfG22kVHGJGx1OERieq5xK9jnwx2d7hoL
LNRz7PafcZXDZ/GE+BQq9fXHDuF112l4qHukNl2XvBTAfGnKY9M+hyi4a/iG18UDZ+xe7Bu05qsr
PelMZEcxq6eZ3lTX1NciQKCj89nYn8SMKQYR2EE1YxSIDKrlnTG+TTKaghc00m7dQO/zWD2vRSLh
J+YcjJr1tjicwOuDI0AM2uleUqj4GCEU+XAccZ/vyzIjzp0xRrJ01eI5Rr/1ov5z5Tz9qr66U3bw
c2QYQCRH5yT8TSnRw3ZXn8VcP/USC3PmzSM47mbcv+TOxMPpWa/fZuoQ6qfder1GV6uZ0IoMH10P
5bo6d74T4/08O0ssEdbhFuqnwrIdKhzXupUFNiz0M9JNxuDzn0TAfwgDRHAPaT9ez/XUKn7GsKZ+
ysi6Ep1m0iTNgwRlh5kWzDdl0TrTWdlQ8GUE/QYzeNsRBLtP89Mhnyvcnbeoakz5lBYlM/PZFDlP
zkq5YHgLwK3EdAMtAYwbIEaDIHXUvUK2FF2K/utQDA+txXzjCWpjVeSksS6pxGeb+n1PA6N1xBV/
1JGPp2YqhkP0p2zOSuVU1WIKcQ7Rlg9MZQMnnUgJFTXQ5CrsvMuS8vrEROKQrqI9HLngxOdH87aH
QYof+xbwTkNPLAp6RdEQ2WZTA9O+GguvJjGFLMPdfjATnyTq8Ga0P/ZUx9EDIWtFmOae3w8ri4wZ
zRpOdiltmj8e6eOz8Gn6firjW6Hy08L/hpF3ONfd4wYH7iDzOzTyvXXkZvALJWgZydfWu7Y3UkiX
LhxrJ3e+k0EVOWOwWQP4LG3HQezE+/3xmYPFFgWv+DjrcfJBpYCKnvCEttODXnpGxrjAoMquQ3N3
qgjsx6nTZ82P7LL7zWGbBpsfyIVIFheiU+fEp42Ci5QQxDbUzqp2sU3ZWW4kx4rGX9EuwsKSJd8q
UpuY4zJZPGssdOR/l+pikpHlfk9yg7A6VG74oD22b5bDu4R7AzfTKdAwFFdZNCu71B9rZCTOcTAJ
7dTu/26XmPAHjiTGMVkYKN/iHsK5A0kbp18xofcJ+mQycs1IyoAeK0DtLhljjJYLgxEjjFsmve+W
2k0Crek/fuWH5IJsZHIFYYXiKp7vJGfbcpJtujIc65CRaukO73eEwnmSqbYctA0kgYQfZBPmgNtx
tJeqPWtRg9xVPnvB6lK9sZAEDjVeysWJ0q4pHpHLCD94vyTb7oBs5qbyU+0dpL4RuXtV3ay9nRb5
PopqlBklCnbt2gCN4q76NYrkWgaGZd4FJsPby7Eg8tsDjvXyCqQ+f5wbbptHpsfaoBZBHU+BZekX
7QUkpPPRPxv9Wm1nmWtbsboDDBhXIRbv79AXKrsjibv0vMpgpBuxyxsSBASEk/yOiqftQIVgP+1S
G1nW99mRi+h/MahYjm3hhcjFE4NHSCUbCNisOnRRARY1Q5Tr6H+BUHv3sCxERw2VV4/Y8V3L0tjO
pJlJGg7RvQjnVuEXPBzsuoHEGsLnHwAIXDn4iaSxIEV3UupqRpTkSowhUiVYJDEmqzRfw3/617x5
aSmXN4A/ed7wdimfsgq13Y3nRN9NXadxUEGToIj0FqzIOZcc3fz0MC0QdN6MT876C2xSvjvOIGdz
cldGrIgT9YDqFfkoyycLuC2iBHhIni+mvoWEXRpiaJDIc47NRG7UbqnZoQaV9QlATHjJ2QPL6Qth
kDMxlVvrLZYU/62cMxTJcy8CQFSAS1s9bp5zAVSTB4Ts2OlK7F5cqm4cGKux66t99VBxmFHaTHn5
qNxwV4Qli4ohwdoPBHBJJx467TbLbvi8QDSWLtaDb1pPUp1d5DUMbuPA3KcHhOQGiM/H2BIGHOz+
ACs8rFTC5Rv67FgdsXVPpvIhsY/5a20qKML+QaBXatRBlmTBFQTGkpa+8Ldra5X8IiP3cQtComzv
aYpsggVPBV/a4LSrCTZszJkhXYeaakDfzVlNspP9dbWPJlc9EDYkDfRJB3HbgQxdKFW7y5MmErcX
q8zIUIygDsf3E8gsOGiERruc3bPJW24IYqZtGfWRGo1eB0qEnbtCqexR+MkO+xi6b6FO95ZDRxZa
gR/wuJN/75/i9KMhynBnpjKRS+CKGYEx7Bc9rjprvSpBdsofBA1D5KRiuh0vUTGqOb5pLlsq3IXH
2TT3RTf01fd7bq3dyyIF3YXZKsM3EDZX+ROxbJKgZa4f2hSK7bS+LCw84de/2epg8OPa0Hr4Or+p
DUZff9+Ul/bnxfP0qrtCjHhTi8BEFuok5wCN0FKsshjFzszt+svtGi6ytA2wqbIO7WmRHm5BTqg5
KtrKQzxPCtNaj3h7/h7E1b/giTr4iXeH6S90YH+ljWjIWQR3h+AexxKH8mdryMdyTeLU+ViSGBSY
haYgl11F9k6sPxne9BoYw030z8vf0um4t7PbfOrKjgwwUggbiRemZIOBqImlFgaSH6fReMznSP8N
I7QuejNNZA7UFQvufyFZDNuS3yn5vUEAusmcqi3vyMa1WLZo0f1f2ZgQqdC07/h9dy9vcAFox4qX
e8idYgRVPESS4VHTxWLIPbOtQP4FLnc+yZREvOPqVTTTxlsfX8pOG4sWpOa5/Mg6WytoLSZGwygK
TgwuLrsBSAcnwEZISghEA/qMELMjDmZNXDjwxoGaNYcHpcYO74lXIdEzPNyFc4iq/CUmYo+svVmW
9CY8pCLgo+RlJodkYPBio3SHo+lnL7wlrUQhUvBfZ3ErP328vmurP4j9zkjqonfpfGw7abCu6Dpn
2Jt7mmIc0ftfol8fuajh/404Iy799xsNsPo4fCt3s3N0g6UCHEi3RlKEXIsEXXpcoYSLCqltn7ZW
oTYtKn0lX3CD1c+arPDaiQ5gUfinJ5WGI0NSwc7Cc7JGli9/n7iObj8I1T5Yaq/V1yLCO5cl+6fs
gWGd2y77/0BEd/3BibkRo4rTgDvGOkKNdRNIKQeKhDyGAGwvCtPb0HMowZBLfPy6QDKdidMQafZf
839uw75/Nq3jV+AgVTm8+LlK55r6mIJZcFQk5HCUtcFbc5VJyyCXWXmHjCXtasaCLd4c2WFelFGx
ytPjtSPcaCTAHuia+j5a2TEBEJp8stzfQQ6Buuozc02Rj1PPmTZlmvzXyGQdQxWURQJDVnfMc/kE
F8oyMb9vqznMGdTMYvJtL2DvuxzHNdcuLlUo8m8SH1llVIekuyHgN8FVLE94DZYC3ep8p3aI+8Ix
eZovK/P1YVQUJy1N0oAfQ40xr7QqkdXKZsKY2W4E+1T23EYjfzhaOri2haN9KdQ5i2Bq1d/613cX
5HxDhhEGqglkPM948G1hgVcpS0fYrI+1zC07YPuueLKlrwb15KFy27q3+jxPmvEWjn6HnulOgFCy
ZiJU8/T7ERq8A83NDTZfoIpKtQO+OnsgcmzYbrfiZ6ESSZHgOEN9xy0OzNQXsjIS0sgdRrFKQDz8
hbA8ulFAGsmj0EaxTuups2UIYvLwVFeIDlmY0068b/rFA/dRo6ycMXLVPt5+R0zBPm7ZXYsrUASt
LUNJ5rSiJXjz1/zwsSHfC1BWhh7G0W1g9hkTQr7f5Q3B3T6xu6rwqEizEE5tECzJEhB5kwrbJsUy
X60PJzngKdLogf11ExLHzazSY2YwakJpXvRdtjB5+ppbZbCGEc9rGBTCQP8BH1CvdnQs2SGZ85K+
xQDmAuEUSdJUyE0p8eXo7Gm+bh93e7e5lqtqalN7MP5TacrlOmHjwb6PUgDF2suXo9mPbCe5VA7b
M2hJXCdPLt6cntOGkv/q5vwUVTMGXCzidgMz0cixTwjNzwgbsFxqMMvp5HKOLkVrRU/RF4W8USXx
LhDKYxfmR3MDPpeI12SWkldl+UudfGrR7JsjMCjBLBwj0flT3PYevI9baR28BJ3VMXuc8L420Wex
47JLEtUDmFkJrpt+aPsUf7tqgkrE4ZNctn4KFOuJNSbwC/i+q9oqIXJeaPhIh/BZq9oVVpooFQwO
LnnrzlHDK4GRpyMEN9dBLLMjFGqLdbBziGHFBcs4tjzblGe881ula+yJT8ToEX1doUnrEqLyLmYL
I6KrPk/DKQlxf6wLXfHD6cJaCp6y1Ax4BMk0Tqr3+aYf9OriObCtxJ5qFD2No2OhrbS+D5sosxpP
y5dQjNmNiWCvGIhIdDN5rsgfLwZKmIw+lpxo4G3+WL/qUuIlq+kIUEy8HEKTGlOwRnizJz14JQtu
u0L3i4ZY2dKAawi4tFYRwohdDrHqSw8iIiFDFk/hx4GOEFMk5F6Qjq2xR471lBb8asSCVYW7gHfn
VVan6L+xCIg1ZzFsi5noFGpJ4Ydt5qTtVJIJ3UBI3Fbjh29MU7cVpHmJKtQQKvrHCNjzRJugk7f3
nDkRSAH1FbOXm0IbdSR4hmPXNz+XU80lvo3qoLTn1JvjhZyZckPM3FNUEzqqA1IHwR0k66uBWHNY
cSPiVrnjNWnuS//NwvXUFKBt/T3jUq1Fi0Z3JFnAqvSweivsX+RtIcub7dgapPBIbIF/n9FFLHoL
8G/Z9TKcJk1q8vhwEUbU78THEeHi0pQHDBibpwgEHqL3wjJ3bxrzly8HNh1rrWNWyzN/aHLHPEnu
r5RBlLCA1SkpkjpvMqnxhaI+FTteP/jdD5XAD9FDTBwpuuL1pIAhjJMo2H55G5UV90+6vtZVYaz5
8QxilY5vgB4qRuDkNZ2YOvNQweyDfKMZIcexQjVjIl8kqEUC80R4/2ClHZWOizfnOrSnjjthseJk
EMQfSZk39wunXq7devMfOc/FRPBqOFPGdYhrFoDXXfu3J8b377pdxoGa5sAHretn5zeicy6ewL3b
MDuWZtMbYLGH8GMjIh1lnDZOVrGxSVLBo047FU+uCN7Q59Kg6blkpLsFuNLFSJaX0ntg/70Rqt6T
mSeSEqoAcD52E4ykjLKgh+jW4fRLCr2YGmCJHrTJffSJuPa7875jZ9ftouE8Q7nJkLhaPVa2bg7P
DGHN87dSiFBp4Wp9Ajcilj1vTnjwVkQmGirqDnLOGf/Zt9o8UXHx5CwoHOGXjOXL1qPeogRZ+9Co
ZP5wUcaIJF/wohYrXteVTbiKR38wL/e3lFOo38GMaMGq/4wfv5sa4PigjLIXf7FywRBGn/8VgN7T
5Ke5rE9Ufq5fHShV3r3TwOjZucZLkDYoCAn+ZE901iJw670CMo2FQZt3UBxwWD3CnKs9Z1vVCgNb
zeDAKBkcuWxVTFdg6rWfAeL1SWuKvmbX5T+o+qZFOu/OTLIrVyA+rzTKO953vXuW9+HPsaRsG2yR
00p3+59sCtsJe6gtuCwViKoiwrz9yH6UGq0UoIcI0XSBqX7mYMNGxm2VgsYlHf1hnX5z++hLKO0p
+xSdcc7nMtdzo73kAvR5Pq7VNDncMxNEkRZ76lB1WVhwBG1Pf0bwf7iy7B1BWLHczfplcjX6lOvo
Rpq09XqetDgnrfIQSJljCR8I04OTFuoWitsZUVLWwmgXBsL7pPaovX4CI6nC+vSn8iaeWbXsPNhO
lw9Eiq9XpdGJF96J8AAiDZGDf6VVS683BztqdmHoojHkbVUsT7x7O8M4L6i/z/rPE0TxxqjI87yD
DNv+2LN5QUk59o7ri+ZTR6JPIXYRdHjYPXyRloqR5QkWA+Up8AW+8ndW2aqZ4GEMnlbCeYZDvnfN
7AEQqI9KCK/hn2t7OHl9CKAlIZlfqDF2SrggtTeMVd5sv2yUcd8AD7pUXBe+Zi2sDsbPuqkYiWB9
r76VgRN+bM+4j5fWSZs+VwONRpF7tlLSQS/Hz/qHJRTZqLlMlyT6NRCmBLqNpRH/ArXJU4lss6xM
Kyd+IhrGcDl0yxUSXKXRnsFTxTxGClWr0ShldfNcTvGzcPGTfSJuSVL4xTNN17O9u4FJOFNzkEWd
wzv8THKtNCQQlyRwpkiLVIeEWCZo68wfuWoZGxjU96l+3pOat+l/QsC29HYvNBwimq/U8+Vk9eE3
llmiSMQLGCIopgivE6vMDcXaudLGBwRzwmxO0gRcWx/mA/Y56uWuxjicvGvhb3QilG88mQqzpG4p
1J2LwbkPwOrf+md9FDYeEXexxLTXFNsnud1Z8LK06KRKvHPTv6Qa1Xc82FLsLupi7ahTSAd6eAER
cVJzhtMCkvQGzoRzldzJSaK2iJvj3eyE15WaLYwB+QFDar7yWdTh8lxGAEPQRk08fMDG8JfrBxSF
oiXEb9elTfS1EjsS/7/plQHdtYb44XZ8rL33gHjSf84te4abnL3TwKpFOOCAsGAYk7MQtH3ThhpJ
038NLlNQQOmi6fm9+e7PT0WMLPTauyLet1CaflOtpt7QCUVMBSRP3+hoXmUYH+t3bpNp/FcsCUDe
P6swr8lZmtn/Ery3zUkg3UPcmD6ChmHzGxhw6BGF5DojS1bqMJ8DZC+de2UX0uNNpWOPrTSmkaPt
P/8veMUMxNxbUb/UwTb6HLEIsabEx9Ix1g0ozONq+x5ZeAWjA/Xls6X5g4KqIZPR/+sh0kJy6FVL
XnFB+1SGCUVDFDT3TSqfCjsyTnXlNM6HoeHbXsHvNS2R+453kse3MGZDJGF0qJaEIcImTrFJKvOc
HNZAdgNaniMdcpVpC/qToOy1H/dBkfypsrHUtkCs7LUc/VaJUleKxlo5A6ZsPo1zYeCrZXj9WC3v
CpHvcuL5K6fvNErluYq2+Vl6E0SpZv78xYlq11ksbSQxD4AeL5+VasNAai9J2QZW5XRPC+zKuBjL
hOhWV6hW4B3JbN8/IKAB5r/jYnlgeujTcorbGTBgaSWKpyw6VVM381uvpYsIzHVHQrRS3j0p/e4J
hlh4tGbK4aiYdobrd7pAXWuGp8NE8gaK/UOf+1mIGUcPI5nqPvJ9xlbEBEf7bkzYj3ccGVUk2COc
KFINa5+T2/q5lFq/hUYW9n3SzbEu5IKUOXs5XcEF0TLDYF7yNLv0vP5L9k0rAJRMTkc9K5NqACoA
yfSiHCAn2Jo9iHjhUtesG01mWvba/uTM41mc19jKFnvkI2FtIDvd3wtLJmEtjZSoXEAfDVit1KVJ
cojJaa5IvYEpZHlhoPVXEf78VzyuS1BeNv5/FhmjPfSWyNESggrBKw6MDhxsj8GTZx0JVQ8G2zKW
IxBXM54Eg/y3WtOCl2P5NRbH0c9ehs8R2drEaljVNQ0kUyPA6E7C5YFU/0mm2uZjgKqXVNylBgkB
yz4Ab2zToBbw0K5NAUjFgC34sUSCNL0C+ekL29dGWXQSUjoo5eK9HtoBg/OvkhAnXekCvoKEq06d
sV1bu+mmMAeBns1u0oEhFT8GDRSvTS9J3I9luPYeHoyOJthlExlw23bqveN8YQFPUF37adxYzhhB
FP4JRCIqW+zGX1YzLhNHmvkA4y/Q0m7465AS75oUhdDXj0mEkTBlFdtFCfzYbOXCemlb7W+viNna
0Pdvluj8stJrrY7tO4P1By1dRpJXrT/xlP8MRGRoSuJfiyzyhGDNaVFy9C7Ad/Iqz0uG6phC1E4v
tAjuGns6EreE1Ds3Sj2BOM8Zs8UZ8lmuiIRFiekPPiV3JmHiGkgwfna0t5wLDwfVQ9TzfO7ivYWx
CfY2BH/5vnDYq8j0S37a1g4RfPSe0PgBaOFSr2zzc4b1xcsXlrdRZFRe+UnIPxB5cg5Gnxs+YDwj
gBwX845cX7raRuBL0nY9+LZhQw37SmOa7468B4i2wJ8NS2pojMmHnVvrTCCyZYM9sdkM38PXB9B6
fqN8tTphTibz8KbPG5AiTeDmeFD3pq0hG6bj7vde4BzCCwen8cOMIIZ9mtn/0wYLxpyvkkdbl7LG
NboRUQBTqrwXAGeD7gSifqIlTREj1Ki6kXvLMSlU8GXuurfX2+QN9mYLwV5KpvRgk9LA9DMzu1iO
6hBdv+n7wdOGoxx3LG1/eIa51Fm5T0y9VgHpOWBZUvG4pEsXlT+RnREAzZIZOZQaXQw/Z9/q4DPj
xuRn922LzQkAGS9YW5h92tftAOGQPsGDieZv6BDuKqAj1TyEnz8EjJ6D2M5KjDn+4RAphwqafNcF
Qqfy4BS+xZ5zRf7gtLkJISkPocDWOn/Nng8hTsxDgdbAPgfB9hr/Ew9VPV9fJm4sWFqG0nHAO/RZ
WS2CcvNSZUzbtB8XhA93
`protect end_protected
