-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
oqtwsV/MTKK+xz+dmnsS6uWbirrIXtpV7+BdL8IaKdksokVdydmYtvL0zzLmNz7i0gtbVHMOpDa4
Ft5FcVYhyN2fZc/wO5b1JXof6Qe9do2JxWwE7iKSiCABdA9n46eTYUt9RvQjvRIChipo22K3Hbpt
qnx0xLyu2To+d+/e96xG+O0bc4Si2A0/Gctd/mNtGdgRblMPodtzKgKkZEtHlzIl39d7eykQYwoV
cv+1hSk6M44EaCDZHiamxpb+n/BoxL4li6l+qOycX4edLNTC0GdeAfRcA8OyOUzWg/Bbvqzgbc0K
e3CLr8SSXiM70str+nb9RKkX4o3KDcy+YXmGiA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7936)
`protect data_block
gblhhh5B6CYtHmJGiRBr13iNOs0TE9PxU7WoS0P3pcy2JX9gBp0f16wB5buAnVKK36+/5qtkaYba
Llc90YTCZQ2X8hy+3hZzerj89twl2m59h0y514g1PEEQi17RamF7h0zVeBWsfMqyoOCZeh+Gl5qw
LuiqVJ1UbGfOyWHxwoxoBIc3kGNrFwbg6+EAcRy+TO9NQ0S0magInRUrNkfcfgvmYRJrguWUh8oF
4ZQ5nfGLrWZqrvcozH+oa9WapDxx3kK2L+/jyYkpMJJ4OQypI5I6bnmyOcr+X2xwTyLbm5I3n23A
7U9hjmH4FSEWuCVhVH0n7mtJEw0l86eJGylLvDGQOiHJMisAWqiVox2zNoPwbVZRp+L9zIRSeZj/
sRJWei4iiZNzd7+ehHyeCD8KTYth8FcKXbLzBEn/ihFNoEjMnp8FjudzujEyZj0zeA4a0A5+YhZ0
Gh6Jh2Ghy4vVzz8Yj86Wa/qe5CvqLrtAhmZjRMIQJKrh2K4MOJHS/E2L5U6Sovl36CNfotA6/I6w
COYWH+hr+j0TCpx2XE+IzimcTN2xewD07eb6xkhlOiUUGshNC8AE7xiD6b2pnPU1f7SiEhWeBgEs
80pyLb1l8HfL/MDm18zjRk8tKEEhseXJVXOengzrgMhDE0f9gXYkbV+Y8aPKQ8rPE5fQpgZKzWuc
V+A0GnxGBLnw0Z/COwJDvT2qsSsaLXPODpdxo3GlduReCPA5X7e6MhFIBCk/unb93vdaPVGEiNDg
J8qx88y4uQNBeGG9t582UPzCtxUcdmXh4HNT1yOdEL9GB+1B7E4NGVY+lMStAFWR0oUN0dmgGF7H
9WSnwlKCX+XQXCLQU41RfIaCs9M8ReIi3jSPbmzsg7VOnkqeJs5vPvwCk/B8qJIXhy4jaTZ/Moov
ergHX+AxI0NsPFxX76H12MkxOL8w+KnQROCfgUQ2fEfmq4XrNjNZlTkJm7WLm9GsmCZluFf5sGoK
tg8K5qHOshGc+uJ54WLHxnBTay6mO73CPbCCzesGu4FyS5+2VYvZpzS+KToFV0F9bOApRXUQPUJu
04n2T0Ui66Mz/uajVM8m688Mhgm1eMhlEYAvj3HOvgmPHS4JH67s0TLZ4rGBi5cf7UmBbas/a8d5
Db0bRUUFjWe/8JsqpOAooZKBxpzQ72EGqHYOzCLVConLk0byajL8QL4XNCpYagbX2QoBrK+E8lye
1LmYjNfQajaft0SMlkHPrRhgafzYPCSlI9YH4APE7IHQlRFCVxQRuZS6KuMNUjC5BazX/kKWE93G
uGs+l3+50oIIBx7KmcndLvGFQFBSsiYlLBBtuxp8iSmqtKSKhUvp5pyM6C6A9IYbzzQCOy5GanWy
tlOn+bCcw/Qp3BnONy+PkuYq1PMuDt/Wz2zmnro0AI1Fge0PH+8NJKyf+LvhaMnHXqcayoFeSE7C
1sU12MQsIBerUMtqjkdoZALe33d20z5im0ZysQEqCu+5q5pENIcP+Ip4sbWnN9ciCE9bvf0jJiYg
V+LqZ7aRiuxKvSFxN/pCFak2dBsUEIe6dBty5p7NtPOXmRf0DW57b0Pk4F+atJHLGXc6r59OpGET
aDbNlOv8nBWhfRAIiOaFJ2lAJIWLv44RHaqba043tKJGBiRHcf5If3h2Io2SWVvqSqLiDxZekTwO
k6NVgka6XpjOxsTJK4BsLpCPCkgh8Y0RgxuTZ1jJ4lbbci9ji65MD+B14clTp03enZ/6JklW3stU
TPr3AwAd+vyuH5N+7l6Rq/g52vEJSm9hUYKIZUt6CEBBLMyZutHO4B9El4LhbUDZ2h+OBX6Jr/7x
HzgpPn4h0ctjd4DSFLXHx14OVchecRAftmQgexZtCc5xxS9BLtEoC+0EGzj6POpxFr7aasErN/6S
UxvNvc065zafsNoK35D4ok0gZcnfFDOoohC2T5nP+He8m3g3I2JwKGI1FeTo43Cd7USY3Fte33zT
e0wp2PPB971nfc3R+UYku5TVw4+JKuOykwIQmEJbCMD3JHqexpICDL4drzw7OA4jmiqQA9eK/aWH
M8UkQX87Qpu7GkYEnGssbQJbGmTCirrZngPAJgbKoV3n3QELcPat0ochT+361rQtrIw9fBQEFaIK
5VqdpzKnGobLDVE50MQ43kTSYFHHY3HaZv0+wm/9vX9eN/CK7DGB85q8wtAUmSjwmokOwFTqv54m
LvkUgDvqXuJRCwZGxjwHgI9MIsc3setqI1swLLXudpRSfhnHLSOUvOExLo3PR9mlqbTlWfgiF1Yg
15iS3fMgTLczFVatTYmsy3yCk10UNUcxOmFTDd8Wg0u4yWypSZXvCTI5DT882yv6pIXMI9YlUxy2
W/DaUPlTmlCYl1wKf0fssOHKDXHTE3HA0YXJ8Oa0JrmqKj0NOvhHatj7s3RLrOC4hteSUXTglfm/
LiJTsPh+Hul9eEY2YdDKWf5iCR1HSYNZiWlpo74l/Hx+5awsqF2v142foc+R3kzT7ydy3kJV+FSe
JddDpM8yLsutR3tX+c1eyUyEO1ug+3y1zdwMdgW77MvFxjBEHIrihYyV52pZ7inVowc8Thh/qHZR
RBA5O8tvtelwJe97Z/R1eDeYvYFkgFQSXS8UPPSFxvVJ9zg0FKl2XF8K6cr+7Gpy9AYgdSfzG0Xh
qHcDseeF2bdSuqAGvcabAZu/e3T9drE4PrMFYA5VutStyxm8x60GCCZkR9IF9/RPv++4NrK1nZLZ
SGgV3ysBTHy1va8H40HvlEO1DN25Ja1PyQHtOTM/NrOOiU5+V9uil3wmGAJbUkF2RlZpJH6z9hwC
iQWc9671xg3JhJS44UvVBkE3Xx44K9Li26chRb6KVBjNcDsllkTLhJcCVF9RrfMpoj6fnHtaaWsE
AMrqCaS+dfYEEgmOSEq4eUzsF1ZbGo0PxAmZoAYYn1S4jM7HBJXCgTXAZzNqk4C5TFWiccYpQOOX
G1+PuLPXym3lcAleHoBW+mPiKG6OPmll079slt1GDUi1c9yhV4A9SSXYQbyp1dH+jtK9TBYmehLm
mCQAYS53JB2PewPO7D5te5uyywjrOxmi9U4VKqZS0nnprt/ypvSA9TyaOkhON8aTZkxm39LE2Guo
nP8hnF9MoVeXWm4fobBMmbn0XgZN7S7z87l4RiKwa4YQdPUmVwdLvbsnlNepPFWTTchmvScniHsX
Q9DgxWghZTK915LqaE+LEMxjeqkMplWOjqsqyVIJS3PShXJbwokGV9X4BFwGCn/jANgdAuvXw/nX
S+y0E8GRulZSh96T7MPgZX2X6+3RxDbYoed2bsm66sSl9n1JPWt5CUnFYDmiwALTe8wSFYcmSJv/
McshJdM7ZGjMEcO3ynjt8NXGQUDtl7J+x3hcUTbZpZLbFUWtjDzBbU33Tg6ztFVNpdpPy/pYTT9M
nwpkLEjwSTB4yDjzrg6Wo0FU6Rvuk6WQLmNTz4v5fVzawRttFyDsMataHMtwXcFzHA4gAr9SYqm2
BXEKZJuhM04M9VJq9UpvY/ATLQ757RLkuNKofvisTb8LRvPv93gMMdonlurWIZyVghG/mr3/wnt1
h300fMfLUdepZaA5S8Yh+9qqNRC/HjND5bKObrBc5GSynC0NG2eVy0dgaK46H8P6Osk5QJubmf7a
HvTMbJf4uq3aw1ohJ8NjsVoCf966QdkVIwVYy200FTLMBNuAEPguQ+KNaddiAEZIcSDSnETq/d8Q
dUc12bnJO3VgCvjgp/XIbIZJs7Hd5fY89CaalBFqDHxEC8Mx6EaVFmBM0ixt1oXFqiDW9c8N6usp
F+KgXzuTbZ/ySfL+zNBQQfGNhMp4cwmvwnnMtMi+73PV1eDyq/CzsoAt/AOEnXaGEYlbkVX1xXSX
xch6yQl8FNiue9/CMfiEjhwjke+axAVGaAUKNtB1kb2AaOlSFj9mZ+w2vy2mrqMEURHcaLftxRc3
TQqs0waD0TGIlxWEvYJiLGTZNncGrBUWJNzSluQDXAHKtlsz0E3ojaLOY865E8ojJFhqIm9f+/3z
8JLL2afWtFH3tYtpZ1yvS65WygXv2mNWcSojU6r/PcK7nYJeG5hN8Cto/AAKyBMZSjXFpO8cIcua
CwBtq/JZqNf19ARINYSZocuRW2mdZXNhCLJb+C7EUIp9bahsT/dmw2QZTrDaNp73lW54uYiVxyID
7EI8h9gb51AoME8XerXHL+DjuAp1XZtIfftdSb8JyFpE8unYleUHMEByYEMlCwQYuyObdct/NADf
E1x0TW8UqqFv5zf/ykIQ0pQ894SCIINfIUXN+vVmJ+jdgInPRQ4uKTg/z9wj3EazRAEO4hj0URku
m2AE3wYnDv/GIv/bf142Y+TFGmZqIDTBfAqkEllsoLHLmwBRR6vMvMR5mzYNsTwEwF4xxwiyilRE
bKg7V2aZ8tcW6NXhYaL8hqts1nTsKRvZ3qCO+MkswYS1lKZ9GuXFcPzqU9akzDlaBchDwAb/W+He
D1NTMGkAcezBz9dXSHLUk8uWB2/5WNjJ5YP47H+DRHWssFLP0RzeEyrPyR/WkiRopMTXVlJ3mtj2
uV8wltWMeyuFtDgicxdJFM00A1cFxY/lS9bWmSX5pQZT8m+z9Rvyw3lZupTZx7mIOjsNgitlpOwx
4f6cgXsaRovdErL/ou2XLHSUM9v5B+alsHjcUGFXfLDN0Xx0XSbwS9+j0dGmfb3yrrkH/sOLcCeP
qh1c2BxmqXrOAPJK+fPogSEasNtkoR4buOOeoZmKolAbKW4VVGbHrR7OYR8TlFj3aCh1i6a3Imaa
T/7AZT/EjuTIrPgNwF1PcyYUb2B9TidqrtH3lESRbs9GaQetVg72R/iPdVZIrj2rlunu0O3c/WbA
6LPtKtvDjGLXwQfNTGusvmo6F9u8lBi1tHkdH13TIRJeJtlsAFOpsA328sXKGl+dATYpesyTe74B
arz5Abs4VwKxI7egU46jwficTWgTkCTpTeMAJWEzAe+ZfaKJSvZM8lg6stL8aW/9uCit6ybVblKe
FGF92tBgeNXPFy8UzO437vF2CYzhETjSIW6uXJ0IqKMLoQ630NedYrxBPCWSzt/AAkdnrpJcH0IL
BFj4l6jAPXzsgJLk4KqGRyUWyKGHzg+fyL4wbW48r7pvZwM7CCmHxAq50lYB3E3jvr+kEQUG+7yQ
q/e9ox/VYBtnQaWyChPhpHFAIsA+wfM3k2UEOsrvpqnee8miRg+C6x6j+ZGXfi5m0BHtXJL4jele
XWPoa7OboOpfkNKpG143UK+vzAQ1vA6+UYUpUIw1Qzm9O885ZlAfRiP8EPhJdjNXjaIDibyU4DEK
4gdR/6vHUOscIdmUStTSnfaVx9m3hiFweGfBv1aV1QdyLwrNP3BzsaLyg+73AqUf9Iundb34W9o7
RUSwKfERMKajKwHTEyvnl7sfNxxTXDsZzyt83An4eN9NbIQm2Bqmu0EFHmz01XEHy/nazjg68Pds
JRbuVV2QRXNIdxomnGg0XpV7yTKlSqNsThzFP79OBxIBzlX1N8r0Ru3MaggYrfzMx5/tHDIF6V8L
5z+TGlR6mACCCr8Bhkgrn8/UleyB3SYUnVsuz2Pn4uNnBMWusF07bmojR14DteZq2bPbWaL3/bV/
uFXil7aWQbBcwcKxbtv+66gqfYLr73QAJhNK+Ra8DSpphS5k32Vcx4Pctyaeb+K7REqfAQP0JCit
E/SuafNnetb3zPpMvmg51m68ZWcMkknZ69PqlT6yROkKjjgfr34zcWwYpYAgEQp/km+O4C98gUuj
jAwcZEDBDU7xvrT2z8V8HbdeQ0kpAxyfaNNhVpG7kfxvgeCoBAq0Wl6rd3TeUjAfm+QypcP5sUcr
XuLUies3Z3oe4g9Rh07VmCfQbgSC5QUjshzXBDNX7ypXhL662uhSpOSfx5RgfSjCGJAuVfU3f/ZE
t1WH2E4mtpkTPdLvdBTXvPqrTOAcVwbLYE2RkroZkAly1DP/yEIC7YzSMCgLQQ05Xw+u+6VfHHmX
q553k/dDD+/jYBDnrDCWS3+KcJLtko4PvY0T4XqOx5dYjWhZPvtiX6+MLhELQJF90SDG4k+PwgZ1
qSScPW5zFpwcH8rg7lAQ9cxR+/KooJDFmxEl7PmeuPOqCp3CCquAfVlS0osf3v/C95m133DM30dJ
jpW8jfjAnID3WH4X3iW7bswXbY3jXYWz8rpQ9gWVIHxhldzDY+DPH6AVG/X2CUuO3J783gYkM2W2
gaXgC5E1HaQ+pgfGiob1LgoV2jUIagjOvK1XvMdFZlG2jrLetJ+dbPQnyTwazCRZygeDlNzf94uQ
/wTHgX74ZWZbawVC2uofnNORl0j5YMHS2xwhl+q7O/CeujXhPjLQhs7Zy98M2UKwpNkXxE6OlymD
aCsjNQoImiUlA/kwG3fuqSjUyEgmhUh9CrR8tWLWpKDiD7i3MTj+w+ZsucuHvvs7cHfd6av74oa/
2Ao0rDdUztkDnWGMMxb/mXTKFkPwkr1dJN+NVEPUqcFxZsZwDLw+diss8qZaKt0TYU/GSMD8gopt
UuarvlWKM19jw2XpbdZwjEJWs3Zp+jf0lJzDpkFiVluEyvxHhb35Wt3rrH7X5AbGGzv0cYoUslj8
9WQeZmcatm8oP4f9SixLsbBa/g8r1uobcZcdo/FObA+IlawcxwZKDeCHd/pNoqB4lWzirl3mv24S
D0q0KNJzMpyOZLssTIE1QymX+3rbWSyJWsyxTvBdSiZl4eBG7GtCEOAknp9+gQHMlhnQO/ERlPdt
/xLhfYOA27ni1VY3xhVt7hJkuGI2ZpwAwMxTWgyfRw4cUW379i6UEDnioy9Z2LKRyV7vgy2YmfwN
0+tyoBjUukf2wJT9kpoL6kWuxLet9FYLtoeEjBrNa/uJvaoj1leaWDE2hQn4y+MyqAJqyuD3zfYN
N3IZkGINfTVoksLFvvT/9IN9RQrO14lt2S1mOGPdG9mAqDx8LtH8VxsT6N3AhZKP1QY0rBz5IsTk
SoHpq7ckhyvGQwUthZR5A16s/7i5pm3V73/P7Behkk5omb+sJ8JD6G40bN1vYIMlmYAQilSo8v00
ls/LdXEi4bHTbLZily2PvZI9xWgJmhaMfCEQQtJSFJKsE2g803C65yg4+FA86dbpgKEXkf0Ky/JN
2mAKpo0/eKINH7aV4WSQgKxJYwTxu4b8NIz3wVX/1W0WyYjNwTZLn61Mc5uHMDGFj2j7VUleE2Ul
t2lsAsBZ5bx766w3Es4b9RIarstqgYWjIgYd3sGi92utYWdbpzfBUKwt7bH8yVsMcurtdlB267Rb
tTViyGMGmnzUjmR+Wu1wkegdRbgoIUlaN/8wLBc//9UwNaze4RFOiA39qL1dvd6cxdngOMu+sJv+
CQYhkZCUp1J+Qdgtl/aPsBM1W8oD1btS0lMWLmChk9pIoOlvpOVRbZ0cR6Q/aCfpju4BrS1k7kfr
t9o6N5N8htpLFSrLi2Fqy8f7zqGt+DfaBC2kjnqQXWdBsvzDejGh/TbxygsSYCjoq3UvtbgyuYM0
Z9BVTLqAYIfE9FP9oP9q+JFyKBRNiT5I93PmOBLdkA9I6RMNn4CRh1qiJ5h60JQp15KSS70r2ln2
H9NuYowqleglVE5qLo+ylWJdyKzrkbdBbqg1f8N5dMLwlZjA6uhNPGE7X/Y6zhhD2F/d/MTHgNKl
gH3J5L90IIPNhHMuMZr1m/cAgoiVRxm1s3EYZcVO8iG8MeFhfThrFQW/pbuGQhC1MQwiXX1Cs84r
fSxpi6m4pz/k2gT08lxqfdcA9LnGbiYICDYtXG8AIIGtNqiwACEuWz903PrQikX6peUwvVVZzYOz
Xp3BG6IG2oIK4FklZ2K0sZzfZcv9YZAkv9mn6J8VEPjofY7obclep6t3VrrWuaB4eSju7s0mAW2L
zyTec6YTOE+JgA8ITvcPR6jihRuVLzePVsCRAu3CoYjBR0p4Rsd9Vk0zmHwizwVT8LT75F5GWJOT
Jc01SS4eFFl2k0pCIEailU2v+2PPjOEdiMF9r8qFOGGdqw47HQu7NolTCq4VPxHb5O10lOcOk8Fd
bB4fjdqwVpizt8WLABFBY0e7tw3GvPEdkfsydcVHd+tRwfkWnK6UjEDoZ1CNgzV34NzpugbmL15t
PcZQxI8/Vv8BKDrAnUNG6PTDb3M1T/nTevsRsHsWL3gTLCRGYxwjpReishHmzkUGGFbOpJfXejdT
mNjuZPsDvEP/Rd9+ZKQOopcg0TbQP7SdG2BPbpmFJrWKTiVbiqbkpF4utVArcPy+I1ud1DgQV86l
8TOhFu46NN63NRypKck/m0DecDVgnngFsgnqX9LpHZzj9qBebPGsym4rgU+1N0ump2+p81rNxgjc
NLM+Rcr043PoQ0J6r3kRcmuZl4deFz/LVIwo0J2I72W6fo/143uN/ny9YWZZb/cd4gHnEIijy5rf
yHuSHAsFGTiicFRnyy6oZOFNYP+YAqWw6qM+2rrRHe87C/iLiDm+t4LJGLR/+9KU1QXXln3yDhpv
foFWlHpzzPhh/RAAKXwCSEppgv/hdFFpX7mNqE662nIkOkrKbEtH5glZAE5fMlspMF9RdshNwLw6
tzPoXE5g5+3aRVUHrAcL/As3bFWAeIe6p64frVb2B5URalwRpzyBEyl4uxDZqOQXCInOdFlS9Vms
FZS6oTgQZa+C+hkGFw6jepeC4zEcZp/fBH43ce4i78bJi1kKY2Cu+KE7GX/M+r5eDU5/5azeC9BD
rqDpnsZgY9afAz8eP8kaEukHV3CucRWr9pNFb5/xrNHmGhIJPxEnM751XQafVWqPTCnGtTHH/21r
o1aM53TWICS4FItsZOYzpr2ev7/GVmiyvpkvGr9+ksW7BGpvcVsWcwWaIKTI0EC6UB2Hczmd/ENe
cR+vVN21VXOmSNAmLC1Z0Z0WN8mc3j2NSTdKigddaym/l8/shEm+Dya7/2BAurfPNR0+bWiT88Kf
yJpKpsn63cOS/lguwQ/4HdcrzmTsKZd5jp9eTdXNxWCuSkwvwKVliXOw8aJ2dJvL9CQ/iW3u2KZC
NK6GyU8AIt7rugEQ5s3NkiJi7iaya740pWGSem8kiQ6VYyddQrqJGFgBmrAWkrtY8RvuYrOGAKko
F3QskLghYWAB1hh2Nxn90jrvMcvmAvRQmzrllhImF+xRBMZip66QwpKeTtCfglIhxSKaW+GZnyPg
37JQutdv35EtOTS8t7Y1ND7FMHZdan+roFQdPscLeyhDwUxtuUTu/tHrLmZKHzZiVyhl98POrht0
AyBMqNcBPogijIJ65ymksRYGep9/k2ertIt4m4vyZA62TzRJav/S0313Al4KUMLFH8ttoOhj6m8N
cVLmAF4II1ATEBGdQa9lWGHFmyCr+XD6EnSrYBDJ/haqZBLb8/R16xCzYxfMBzTxB0XIuUFLf76m
J1F/NqJLCnRBF37/C72xSXqSV52sdz8L9CNqTPXyRLzJOjm2fawzuj5jIHTzVyRTifsG6ZRdM7lb
CfXEfogM/whTLMna/IaG3scR+ja34NT90kOgkGcwAdZEO9qAvSMtnHRnVuFoENWx/NM75TLGE6km
n+1+K5zV31+A22SMlQqR4ktBCGIqJM61RYLa9pLZfYi0rGPSyLhXHN75aVsJYrZLh6eUm0DtPFnK
CIwaQ5Dxo2W8JMbU0BtUt/ixpHuIsxQ/gJlMw7rX8q1t7AheffJH0d68ft/7ZUjelgCDG1RVa7bL
D1EdV9IDGojF0h+pwpEtZzkdbMd9+sRJIPfRDors+m1QRwImsRr5z2WnBJs33OQLcotaJA0NCwol
EolYix9pyt623/3ImY5gh+YhMrH/PTZgXzdxwRZgbqKr/M2S2Lcyo02FfxuCgnA+Xr9oTLvJlugz
L/f9AJ5CibLpKuUogkbbYPn2Byt09CSfOKN2mkyOz624EYMLWhMLwKDWMOIRCeaR0GQvOvXFk9PP
E1eJ/dT1Csuban9W/lNSgerzrtCBwmq4E98DIPeCZkUW6A3rxJsKu8ViTw6xgJ4WK1fIYjliCUIc
RJUm/B9wNs91Pp1+6uzzwAF9v8DYDxfurK5FAEkYzhCKo1kET0rVdvzqVI0mlJIU0RK2SngxDBEh
TVCzOTgQZjyXQ30k2Gj6XQLSaluBp/WUs67wktAfQvhR2wZEx5GTYE/xiCXbihIkjVsms3y6AhEl
ioUX9gzWifaaxGzED+rZBs7p288JkZHvMGAaNLCV6bSkzv9akF+PuwG85cG1h3OagxjKkxh6gxYl
hA8I8zkQwLzLeGdOJMg52H87kSqkG5gPGUVnb5dJ8BHX3EhWjQfJ891wUF3dTaWRPJzN3/Ayyizu
rmfVLEmRjtuvH6/bTl8VZk/ze8dqCl1byLxuWrMzD6SPgOICSo3dR03/lhhCxI8vOilvzH0hZ+9j
OgZARg/T03b52v9H18hu1kSlk0hXNcwGVnIIRYSV3spf+uRXlqHwrjMl/4VZlxETvmPBkjyHuiPc
NItUfBqk7PBKktyAtkJYP7D4YsTULfIkAMhZDC2nPyL/ESHqO1PiCikuISMEPAjehXErRe3RslB7
FKfTHc2wYw7BJC8srg==
`protect end_protected
