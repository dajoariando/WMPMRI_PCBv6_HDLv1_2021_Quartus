-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
WJgHnTYstK8IkmtFS729GjUFWL9SVhdbnvVKYuCno2IMziM/ctkXZsGhzzV/0dH+SwH9xi52/BXR
Uh04yiwhhQ93Dc6gUKAh5l6cu/CldGqhl2BT1VyonxDaR3Q2Ar8lJbJ9JqQxFmyrgDnISuvgfbtt
l3v1ymCfpZNEudZihhnfmwgTlM9pHxy7gCKiPUPfHV983N3pIi2/mdP8Pg/wm1xfMoVnp+KyzQ8U
CWB9UauGQlWod0r3YTlpexUbNZkbrIxQBVeZ4E1XZcMtyigUTXJWTRSFfNbqywXow4EkXlrjLHPv
+G5koZKro0JXPd5EaG2RYjqJKrG0b09kEm6X0A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 35616)
`protect data_block
MeOWVMhyiYaIlvAO7cStHdFtCeXiims1pvxJZRqfZgB+EnjKps1liW8LWSiPNa9P380vmzsvyaiY
Y9xLixgXAi5StbQA5y74VtQjZ7ywoWhrLC+3c3MzbmHxv0gA4j/+rryRQx9Mr6W9ALwMuL4b1uUJ
mcf3ONO+WCZT3Qx95MPm5jfnoVRl0ikrCzJ33241/ogoQ3Z1wmyCBGl3JU50hM/udsBtMjp5aS+N
9O08KyyFyzrkvdSYWNN7ZKAxrO0r1S6nvme+1CPMlqGmxgW+/rVYLrGNhyR9urOB7N2KduO46ID7
CNWdFbJmBTLw/z9ugXr9LoegDl+sgEEk2tHYQTBlNfWEc5aw+Ls2fZLWSJVwzvCvS1WNGSUVJaYX
L5zpHfQ9BYqxunFRNnyS8qEHozoVlZNzJ4pbkidGTP8X4y/N7L6Ir4QfLsAdnrWL05PTBTtFzHfD
TxzXn9iO6BoTgPKIHdoel76nleGzfj5xSQnr8axAH9lJFCykruLG/q81Risiqcmd8uUBEIBaO7c+
HY80+51uhVuzyu8//VRaN/aETluT4U0pkWzYi8yy6cQ7BV0dBtonRdZzDsjFH5U99N1qy7BHWzbR
AErvP/+uRWj8cofUMXSMsqsXnv/b5jTB4sbkvX4Y3c6JGJ2/fbG0AcmQwCgfsQD8rTMr+Mtyp8bK
rnqhZ54NMUKDJB2Ye2SjSWs30alTHKFoTEHIgaEj8EWJrWK/OcxMmzKqXGftEbF1vQC9aeaw0Rs8
3pzQkNHyvvB2qA/xdhGgcKCXzpE3bcS13sw5nxpMpbZ8IQgfokNUN9IbRuvX4yTUYyvf/Yd9QPrV
5Kc21M0mIZCUc13JPvqO3QyleHdKtV6LKyvP35d3NW/CwfG6MMtsxC1fhAt9dS/fQb0vSdPznX2l
kUuJvzojMKtVi9qApzUYk6YMZ6dkKfPG8OQsnpSrVUnI8RRSsCHgVkLyDRIxl6g4UgeQOg7atROu
jXdleiGMLTDO8cWthfi4LwUIakxz8xQQNmSmGIsCKit67ayF2lhPkDWfeaOZPL5CfYL39G4fXNLc
aopd0/nBLXSYQvmIimAfpD38913nJpzcZsdA9wyd9l7dvB3OPgJZkZ+9FB21TKpmiSKu8iRonZQw
njQPi7Ai9IzuiAh9aYgGn1Vfw69yzDsi/HCh6MDOmTvF10ELv51cbFzKvs6pYuUaNfOD/slJyZY1
cDQfk7H7OHG9VLUMOKAENz5oFh1r+zj5sGeUGNPzR/Zztl9Br8W1+rer9rp6lhQtrufytSZDUPwJ
i4YGqcrohTBqJGSw5j2yMfvnUDyL5FareSZqHr91x/lYms3Fau9BUG8NfC9Up9B/McupqHfcl6w6
nH9fU7QKXEfpoF+qY/vDYNvFy+jd4yGZCSGnJcrJGNqy6wWYexSA9lQDjwP9S2JPp8E+y0qKt+aj
IH1b7YnzYIHi6dyT3Vujql6yu6WLI2l1WL4Ogn/Q0byUOfcvgHrlLXcDmw/MCN7gOrt27NBpHUC/
JvccPPj/AdZR/6K7GTpsUF7WsBzBU+L9JwMXmhyu6x1uzVSQo9vJMgPqeSm8otoXq5eG1Tf+EnFw
+H9IYPTaTcyZKtv2oZTm6OV8OWDpDq5Dm+cS99jT5XUmQrqAkrXQzL2xi+GrcXxUM/jB304++i57
wbl0ZQAweCEsv0gGbqw1+t7isAsFIIOS/eHTB9T0n/Nxz7cEuqiDhy+0O7VK2njLFw6/Gy4vFZyD
zQySTPE8LGNdJ8hz3SkRGrK9gS1mG589wOLSLFr/UgevQprHR8Q6iqRbDlA50580mlSItA5BYLE3
uKyyEhuiSNV9Oy+9HewsnZ3zESWUH+2LZ6iJQy6JSfV7Y1asIux28G6GqJTK721JTTdt74/rU6q0
KXObAZkXxRNG+4PRcXi0QzXqJR1McLSFJlf8lHaznAsyKsrE74oVC80dLOMPwJ1Nm1wPwYFjEBcS
P+ZKa6Qb5s0cy9dMeMJk8XifJaGu8kLRuNBOqvRZGcLy7b/ageMBiHbBHddfWUDABTew5hxAfscZ
z/G8eQ58S1/KcsomkumsQPoiFGhixLM0ErbJFb0I7/tY7kCNbfkaCkz1xoB4SVbwxXI0Y3otYFiP
ueZz9guNi9tgskwUkJTFegPkCMjoBHOn7Cmb0dCwd/K4cosrcYsTmJZEGm82Aye9e/0JBtVILBMX
5NmHF2UDlftgPqtAEb0d0WPexShhZPLJ2QzaBMGam1DAmh0REU9ux6sxcalelAsGPxIP1Ts+efEr
SDcgG7gDr54O72obS/GLIj7Yvq2nOMJTN+fRBzZ/yzbPlX4U4oj+KxtxHcRMmWdEZQ/jiMKknVSv
JBjaD/rywJJNBVdaChkUBJ4M0IDxuEDhjU34x1fQ4tqrDlGfUK0yQs2NUkwbwuGE4OXKZWXnGPfT
1Bw3w8V0mZUGuiAQLkyD/VX6irEOj+Sdmj+zvc062T++RzxFf0hh9SYFphGRpeF1leBUC0vYJv1/
F2Ln3UQQa8k+jmCwRVPb4DY4zc/eGF/oSkp2wtYLLPjfUSIR6kPCiuLC9tFITmoaFQH1fHAUZ7if
V4u6D9sMyVCpqZ1GgIQk8WLUDj4oQq4pe7MVQFGBSSqY5F2Nxhj5wFBt3y5NcfT39uYnLuFU2swY
9i8McbXOsW0ixOeq6qvGDcAo8YZRGOrKiLVKq4wX4glKpkA+dQU5+/pVw3Lrx7OzxV8FcYMzOeYA
CD/V6sDol9MG1NNrv6vLJ7eOMU6+Qdl5rygedkU36qPU9xBQPPt2IrAqLjPm2qCaed1VTRAC/8Bd
TEzc69+sCNFyhrEZQ8E//6hykvSdkKBF+ghUghkV3GzUj3I+DuGkyZtzKilnffZpr80DySPKMMcf
+MkTsELH2dp0z4dFFXvGDWrPg/7wOVizZ2rGk1NIRZ12QXa8nVCc5h8Z6G4wm8mI1F1k4wJ2IT45
CU3OGxh94j3ZOtd9ZdS40szR3zcWzsFM76L5u5HEsCy9soOheuRxY3oUGsdohviEwHW0dngLDWrI
vybf4bieTENnXwV0kQ6fpEPzhWz2HJub+CFQCzXsXwvLoNHRvWg7LRE8DKp7QPt6W9m+E1ZBmulq
dGCdxj0lnySrTQAlz2O1ottxdtYoBHidsMmD5LVlVsfy/0nwn5DbCCvXevRfYfYBNAsPp065fAJ9
6w8rku9VXxX5W3HWVf+FVqhz6hM3aYVm7UGKtMZaQTXDp0kzs9MxaoRR1tX/TbxCxN3U7wFcEstw
UtVI9GXIlOfpOmSeT3uQ6ld0XtKEROSDkxmiEOj4pD4FOShLFo2Fku/2clDeniYxM/uhFFWhR2zn
oHPesfxpGteI23p2Dakoi0FMD818L8u0rW5y/uzHEcUuKyi7CrcYv4F3JlmuLJKXpcdMJ4jTQxMg
QXsc+1edTcRjPGLv/EdgmF6F3a2vcfWOmYCKbe710R5u2Rupv7JlUuv2NyTKfbgrWlf3IU1bcta6
/rhccXeu0BBmPXXOorAQVsKTmvuNGm3gKESuazclC3f0kyf+PTSYdLOh+xoEJ4TGyiXCZxxyxBA4
xU/OeTLLFwGj5J7PLryypTi77il438635yL2rNgt5AQeg9JGJ12SbQXTzKCYBHbro32v2HXWq5D7
Q4fv0OvJDt0582XFDJN5L7GVJ9tIxCHO3HnISV2ct1iz+K/oOXIBtjdPK6y0Rqmj4JJecvuQ2JsC
yiJQ5xjjRG/BV8JPlVbEJUhv5EStuvTRHCqT1ipOv3LVuZcUUdQiA5otRwoWJVyTYyp6he0Kl38A
21eMJN2DZaZB0InGd4iQFHwL+mMY6uDocpWypL1AMbb5lDkLkcPffjTlPFjpV9Fbfpu/PpZ1H6KG
wHC5bqKtNGlGWceGSij+uNtmPW/K4kL9B6TWqf9xdyWvNTnbtg09GDObrz8/ewrp8PwNp4gYoffv
Tpvb3RZtX7njOxe4IXtjvGu8ZdneWgdcwvnczGEZ289uHB4sSyrIImrdISy029fSMAaFPvL7aAX0
T16JRLDhDQnjS5HQYP9xi8TQ3UsFPAapFz+JnXeutmk8rrtVWaPlNHpciWEH/rsNfcIqnfftrbI3
v4oiuv8PZ32mmMS/OTFTrkSBNcnThlxerGu8fCmWJ3bY2RSyCWq0Jd6b4eqso44unIs08wb/5JJz
gr6kNJpQVBwydfcwI5psrXONXVLMYBewQmTUAq2NRlusKt3ymSnFo/UW2//I9WA9P3813E0FyeiR
z8WVF85W643DvUq3xy7L2hsFiA1QwI9k2qqUuYQ/6O26axB5TSvSEU27zbfpR933MWJO5OPIoRao
0VUDRUYbQwbpDN4SWewJcnbQIHLsBNBywgnEHLROpBdIyepi4uI7nxPu2HNRUmKHudSVJOJFMRfo
F2VPxZd4rbaCktza4CSbx/GBBOpJrI35/hIXmijGoKs4gklLHncLGTi1OQykCjqspRjyiXUConbP
DRrLUhRyXX1Fyf0Ph/BoVlnheRdLVG3BKrA4kiEDOVfd/UqzXjpn+6ois+XajQxKSnEjINxyESYO
lk5B4PccKSouEaeAbkkNLptaaBcYnolFWJ00DIN9yBKRmYMEN8eVQkSfBVvyXrGXMS3dW9Bxe0E/
RMkdArGp5QWj6JnG8GKj+yQ72KAY5h7MsGH/rlVr3AQeBiczEt2r42AH1J1JNlbFY3JQes4XraVS
PiuZLvgl9dTqFDDfAGGeyfvXhWg9SeiT9cVTdo5x0wcG04z/zCdCJswo2aElAB3Llv0ClVUOtXBM
hyeYyOMS1B8Ex7jobscGWuXOxZUZ93p00MJyFVufRL5k8Rx3uRTF9UAo8QnQYIHWtEzDihGWNdoR
hgWFiCBNH9bIoTLpYg3MU4GSe6ssseXPSJZHxicVbA5h/1IjKdTR/ae7dy5ToHuAybIT+ipmsbz4
bVdCsIRWl67Ox+yT+bYU2Ldn+3mDqY92wZrham48kq67za+f8W1HMo2NbCCagwf0fQPNTrXmbLbG
Q3fY/hEdU+w2vTbVLR0jI0d59JMIEYFz40S4kZCAAL+evVDvx4kz1FnCozUa50njuMl37imFwNfj
WZ8CovH4/LNGVmcQRArK7ME8x+LOKNi0KxM2S+G7aLTNXY23S6UQtju59hC8ijXw2nHVWvN1zD1U
kZ7ay8uRkaKNMqSmPFaateeoHX5HbEtfUONsD/18kNkiQ03OU9AXYds/oThA5ZBhxNJPysdtKnkQ
MbsplDcn3MZbHjdgnMgE1lk+nyQcvc6GuWwm78VxWhbND+zNhmaBcNKxQpNSBSsfKbK/N9efUUIe
+iD+Muukl102BHt5HD6xMH2bQBvEEMRXkoAONhSzD6JIT2eeWsHgYhgcDbnJ0hvtPunaBzCOlOU0
WHzt4c/iLEHHaK9xGVaBiIvrp9mgWP8zgYk7RJb9Lr37so4FEWEMjuArAumLKlEDAFNn1AxDrVPp
sC8BJhLdMC1lg1Rx9kGTrYakz3PfXM3RMOpw1p/Qg+R0SGpRkfcpAWEJ4lgNQojHkAd7xsQg5VOr
v/nOOneB32FDXIMi+iZjQHoqTAMXazJGXqqL5JdCxm+ovwcUEE6DaRFcuKw31OdBYttoimnJg9ni
hkbqtfjscrGs+EV5aDQAb2n1GqCwkEcEuyFrA5OrZOwJh7caoq8j2oKkrME24sZi7J/bbSwGOmNa
eJBY3C4w7lrKwlpZ8OEoYy6vfqBobMIlmJ+W/u6Jpl7xY+30FKWeIcDbmpk/gvxm6OmEI5+rSIJC
FfFqPtOZ1sdoQEYm8vr7gTQpaOIVKDz8K95T+qV6M8yWTeVSYOEhoxPwOhBT5zU+4RGUL+1B9Vx0
Bm+INSa+IpU24NWW/tT7F9Sm9ePgkp6zJ7/MdM5/DK85+pOQbVQvgTOQ53q3LIWQLuC9qlWqv0Hu
/ufSmNorKVwYrsHmVp1xx9QtiL9HUiDHRdnbZDl3fouZANTi1dSwcXxObRPZuzTKItg+JknZOgMs
crb13G6phRSeYwZ+/nNbRxLUUmQNv7WXudCKB0ZTgDPxHHFGOKQAt3EV+ffsagmhFrCi95Cv5lFP
ilhd1sP1vGWlAf9p/TV9rXQos7kh7cLWX+wnN0ifNTlH9zozmbtsEjhLVQf4i8Dq9wWK7++9KR+z
BzTnqRBYH8tgrlCp9o32GZuqjCEyE2q+fptHYuXhqx4tSIGj0s0GRCI2wMhHDd+pT50uPTMejmta
BPflUZP4aIPgyYLQpMnXEcGjSkirLtKdZIL1QLg81UDts+tsqAjDmMNwYMUGfibod7tEIEQUBE6O
ywrhcDqroO7r3kE1oIfxRa3ewMiBqZj7SzsFSrqXOdwNuAUuO+ZVVpDgNoR7ufrWZo69aQLjl5Rp
Z2B4sgwTJVtf/AbUzARhnWJj2JMrHQFQe8diWs9zvWuqGxWoKUAoI3TNDVsfMxSFOmNwdYKH6W6G
NbDSzBDZ7xV+HB43UJlybVTVgvMHw9d5Ulz0W+X6CETnxr/7l2dJJqJFZ4Qymc35pKkIGVRQt9um
zx1YPqJN4UQWY6D0NDRg7mK8Xo24MlPdqah8Sbg/I7zwYtD37rOQ+3fbXtJGHJe5FbtIUtw6+WJc
rTH80N+HSSsrpDLC/XpiVM8fZ6XP3oJsvSrQs2AT3IiE2vEMW6VISYYwSBkegeQ6ESG/mmygKCM1
VUiYmgsdBfNwOse+qglJ3uyX8aPAQvU2TxoMED3Yi/+WKfKHNRNWrqTM+1V/+MoalTaddHDG6A4q
J/tGyt+I3Rd9Vj5sg4M5zyar4w/woDENefwB+f2UwJY/0pzEBybZ6so2a6YrLGfuTn0hD2OeJSpp
txVdNyK9RYNXceuZM6QvRBxChRT+K6CyprwBMUAiCBjh/+VrYNA+wteRsijr6/gfhxir7zaaGq7Y
tNQgPS6hx2VG/B1XiOAg2DzEJRiYSvYhtVNZq+Q5pUsvOVyisIHdyiztE7k6qnp4Ia+zkTrtMOdq
UBUu+MMbvU47qoJgop+QG1j+psum1poXY6m6mU/8T+znwgLsP2nWXMBsZJm0WAJQ1YbPyoSHndnL
e03cuulGPU1k/4dvs5uZI7YfncHLcnPlRAkvBiNWC4wlVspM1RshlVoJeEhZpf+ogjb8nDFvlyWN
JZQ/YHIOwsS1sZpY03nFdHguFuckw3QE+orK9O40Gz9GpJu9V2ayFO9Ts9YLUgYGZCDlXU6mm/+w
xFtQg3dNorjJ8AyA9h5yPqFubHKGl59d4oPjX2+1BJKa5bRUFGKhGP9fiCUaC6zZ9fVcAIeTe7Ws
jATpZz7VEcNLS0c143gt8XLmWW6ICrH0VhCtDmv8e2H2jaAvdtUtljF/3bGSHjdYLwJGyzeIqtl6
u6hzPpMNPyjXuNYNrNC0ztrqBKfLBJn283JmGGxtEaJ4Jf6GObP4d93oX69BfOOdbeN59iNre5rJ
tEvsMeuycqCaTiShiWw5jzDiO4AoQWJG5xMjaKrjeItE9oOtM7jS7vrVFHvdyDE0m7qXlhdpFLSK
T2nOOaAQGgL9L1Z6Mc7DBQ55cjx15ROjeNosfVzkJkaOS5q/zlLslULv8gBrlhUziqKjcjJx+YNH
ALCieWuESye1/PZWtXTBVqBrsblOhZvimfn2BrhU4QfCYoe/2Z+0kMW9PODkBk9TTbNGeui2pXHb
nzhmQyrX5K8oeqcUDwNllpwb2NaPb+yi2oBEWaG7HzzAsL4elDjRDDQ84YaxFK7vk750umESI9W5
EHc+fvdMxxsvlYoA/rbme/ER3oaZuPShBQ0/NBV3pWtp+PMb2p907ATg9IY1Y+voZF17RX1BUyVV
PzdDH7NEskzh3OsGWk9hY8k//ZOc8lwyZo1cZ+FKafKGGcbQcWiAVSTtu3wlsRd4YGElTJn7G+os
hzVPoXKlTfNiBSVSszBYTnEBSZh6lw4pnjwbuviWsIMhccWEDv6vh3pMBOEGt49C+IKxFf0taZN3
gNMw/hcqePgeqQifP+Q+vdU4bFZF2smcGnQCUKeWXvHqXj9sIotIhaxxCiolI4cBIqaiEbmz16pJ
f+T7tswORSse1A7FeT+gifQcx1aD6WmaAbNeM6LPOKqg51AtDGpBZ0Ioax7K9SQ4SCcF2MxOnT73
SfwzSXw8zrumupOV+lhXJ72WZzCYlUJX8+C0sSTIwjiD5il+3W4c3dZ75etvBh7JmL12T+PdHvzj
8/JOr0YnwJwj1nHnnHz7OMBJvMQGSEdLbU6JSdWjYfs8gOY/hlEIiN41vx3HeCxvK5SRF7G7bPDw
MyNTCgSiToOaudCO/IU8ZVQ4VWStbNCgyZ9W9N2mcXN3uRfSYGMFafmDmJTk+klAkfDhW+D50PMU
Ioi9bua1IshHXP7zrkT8OzIEetWVJW+6W6RJdOPNAGrMhmarMPAz+VdtsyptGf3D0i7lXH1QbFTy
m4OFcLRKTiBQ/OIYPEwtepEcIHnUJQZ3viLjSqdropYU7rsmzjzKuDs2o4///3nimVKYgYJ2SZ8A
I7njoXjJbgo/5FiHz+NAiZ7mMV79ouj81OO5aClawNI01q+eL2y5W0pZCph14yigpHbtprohpqR7
lFf4toLHmNDuWps+fi+nlK3P7wxNEymrET+V3i9KwKHRHclXxEVJLJ27XnCkhXk2N9FgzbBKxu4W
9QMV5Qhl0E7sySbBPWva+kMiF4Oq1Mq+b389Dbuerl04Hob1szF95+fArAxB8FCGO6NefIH+Q2QT
sRBtgDVSbevV04bnDryp3FkZacOKHo+kxwUyWYGI8elvR9mbYodhQcZpFxsNYh4/G4N1gVwpq0ST
8S76gkwNRRDNP1X1wmJQeXFOAHElCe0BdzSSwCLcwS60RWeO7RbKiOJduZi/KkuRC34U8zkbj/Yr
kWOelRTJ+bhCDqYwkEdl9jnwWf08cIlXOJzIfs/G0ojaQyaklml/pslxNIuh9UmmBt01lcSjHVmQ
GzANg9kEu709yPCGgAwWZ4NsARSK++8PO6W07PU0vkoaUZgwRAcU/fzPyh52okcxWN7572WKiT1K
gSJJKL+B4ccmIFT97Ab4uzVVlbaHDeeuqyqIkQlCgThYKn5yd+TYybqKxqTkwmR5/vGsoRCSJocs
w6ew55rAgYtvJ0bTjmTZ0jGu8l5sgyHbM11RJZJAaj6nbV6yaveZAD5cDu87KHi9PFL92FCCRByq
/+G/cwnfZCJBJwGmxCELlWeZbB5SUH7GTuLacRXXFrV26jE3gOkLjTyvOQqWfPpDDRDlHibmQH38
8TevyJWJhWVRYu08PyrNH1AM44tT7SEwfDeYMu6zHh2Y7akk/tllWyV4bTZhe9gGFEa+i8oP5DqX
H2Bq+9YRqLKmb0IfJRLQE3rA/9KlgAqh3YkX6ZgH9BLKs86HFRLm2RhcBP4azSRKQFE6HmK0Tm+i
HTPFnRIY/Np9mVzDcUWOCBVcJQtO72qn1KITeioEIb7qDT0YwoDtCAiHQvW4P3TqzD/2DlT6SLrP
okCGamhWV01kVUMV3Ha8ppwSwli/MldJ/GOtxxRkjx8i2+Y/5W9wGyOEbMBiVcsiwazkcwaOSdcd
2fOsLRcvnsfGlODc6wwO1EHXrprpHYiLqVmoW8OdqfD8K8so1z9ytcL6Jq1XDL5vExic2MEXRfL1
D+7xObYpyHWu/8pDJDWwS3kOPIyLYYFbs1ZoqUZQu5lwXmU8ktz3NtHme9eQHu6XG/cH6ohgGd0K
w5WurhLh6Wal76EHh63t458s1u/JbyCKHi7vL1XuWKPcxk6n7DVAIL7ERNoHMcME9l6KHST7aM+q
MGDNEukVzUrsf+6v901y2KY73N40BjR2XDYfqKK6Q3EktMvs1Cx4bjPi9ReXxSgp4uLlSa+8Z9f+
k2imaafbbEId54o+1wrDrFAuZJm/XrsTPbLaeIlHcHWw0eVOiWUBwrpudcgVByZ2grwWWvyCWix/
vnkGGbkmgFMs7lbjLxVMANAGLvjefA4hOtMCZj2q4ZcgE77WFo+K1JL1TM1gwYYfFzWQGbeFLoyq
B/mBydQjLUXDVZb+NZiEI3D4gSIGv03sRYNB3ZQ3V/Zy/RQDPgmjV9xQ+MfMV4Qx4BWpLqmNm8KI
waqYiBul35HWuCdkJEn+ncmC0zzR2Y4yZUI/0rL9vbxUjM7xJgbXJwnNxfF3jfkuPmKvYts1iJKF
KWazy1uOQlT6WZ192QMcGowOw/mid7cAvAXuh8TekPHeDdWaVjNdskaCW2ykZ6zIe/fKabOtv0UT
nv/L4BIJrwIMgamZPYyq/JupVVIBHwgZ4NqXKZwqCsTcjilap3TXb1/OYCiOreRfa/3e8JdBkL80
yegAmVw/HFWl+6pNxkeDXxRp3W5djJ+1bu2r8c6SAPxb39ZgFwqTwV05SQPNXgOUOx7gq6v/PkA0
m3QfWzXonuvZmSUQOWiv4c4/hEO+JGJMU9SHOUbbBFsmkoLLdpg3CSNyLkIV8q7UTfAKp3tMT1/e
A+5QujnJ5ZAQInzDztqRcOLjp7ejLtm4Bi2Br/eAnmop2Q5VgAspUU+9HmDgUFG8VGpBV/qScYOB
Le4N+UNk+lm9pFGK3zXJKpAy/vv4gY8JNHnoM4jsW788oCAKhLBcVETnNIMRACDSsb6JxSLdxizm
FwQUWr9v8FCb4Vj4rDb5NSbuV0ML3F/y8TkwDxLhxxAkLPA//vUdqTTwb/XBWBQiJniFiAWx+P/0
BIxmdgBnIsNaFuaqFh1Q+oHF/iRvY1Llr5qZr/9l3tPQELdxJYw/HrcthKHsLbSGGRFUZbRHzNDB
8cr0Mousl/F9HqZzgLpWXkOQde8mDnPfjKDJzUKc3w6WcVb/PFgmTC+SNiwZxRJKEAcHpP6kTKBy
3btLrh5DjMsIXgqHmdRaE0cjcwuL70Vfug4IfSUAetm+ctv8F7vQiTdEu9A4izSzmuDXguyLkMIB
n//SQVsif4iWbR8vCPmwBJWDyyHHSdjfcJEjw069yp14kZil4ZX85xxprQDiDSo7+8QKNXZ03BE5
MqDtIIPsUU1r6UDvS7N0l1RqgYhoSiQOhbRZmj+x1yOGcwJvvl25j5toA4Pn8EAnzrhV6JqjaB4T
rpu1aj2a5xxbjwSUgUd0iUPU/zf5Gztba5P+Vb4slYf2+q0DjJ7mU3DA/Yv0t6Pohl6szGrTmsw0
gmI01unFl5H6Rx9m0Q/WjRSeisJFEhrvCa13EZVLUiQFRM8WB7TQO1aPG2692Kf9Dfl0QqumgsYX
+cRb4pTYsIjNay+0nqS2rqIpk/Q7oOKbF/wPkAy2yZLOQFI8SoMe27wAiK7iw6g29TySMRhEPIlZ
BH0ZprGz8C/8/HDRi8wkwXe1+WF3HsZdyQ6STkiu71OBBRZb3d9h4T+QwvbSvsvEalmhZxhBwgHG
nCCNF7w3HlDZ5gCQOBSKq0BQNJD6HuWWkQ6GO/73a7hJ5qi2EdK8iUsNWBdUZV2KXUo96dH0EkZp
yF65S1llZJRaadZJQCRhZyBhX5W9nsMadU5MliI/YwJgeDN5T/DCrsHznGKx3/b09de1H4wHOs0y
xG8L42NBw5yAD/46na6KFnXeM6jmaVds005FdgjHjyIMPmhycKfU74I/9eAAs0ipnmIWFYBXok6+
FktpH8ltHTyZG9zIGQE8jXQgOclhaLWJhzmtZYH6c9ky3lIUMsSW+yLIjZQxtG5nODsQU1qlIbIK
eDXUOmaylFFUrn+FAksXmH8S7fZsJWw64NQgZDYOr5aQscfH/7rdLCfQ7kP5o9YKyt0zddUxRn6Y
uqWbTbX0qK8eQBpZ3tXB6BXcIiIBEfLC0drGAxyvqtGNEV2R/6jW+3EA+HQq9wAxrtN3+xRQYkik
6XUulrFG0FtDpBIChel8BcslEAYHHPeV1QRMHAFH6kqpq4uhunKiSYFJMCOMc7298zcHPmVrohKk
8Njy8fCvebDPds6fg7hMVyDJ4v1MDHWAYXPCWgq9mkrsJVyX4ILc2YkIzy59bLH+SDXOJGWYM/9Y
Qj15tJFOm/aC3BTgwlKuJ6BDFxlOzBvZnwGqyvMTZs+NrO6cc2NOrdKxvXgy1nZGphvWRuYvwkfx
N8AjpjwM8GNztM9L8Yi/hT2NGoiR9kGhU2GFwLcnIC2tzC+jnDA/k9StxKsEUaBuyoeGV+AksXw4
Q/l6bc2i/3loz3xHevHnOkb7DmROsQksQfi+4Q8iJYqXrMtDK7ZLRN3Gf3nN51PVQE/ZYYx38BKZ
cQ1XWMtnekwEeFSS+P+1I/m+SwzFjycSuPlu0ViuXZkTNGWrByK2USJIwx+sMXVAGQ/c+m6NL+Fa
iQ/4a7etM61KE/CDCqcFityxrRa/K0SwA6QuDCxy5L7lCP+KV01L12shSQlO7VrA/5nHJ/BFYvaj
M6KnzY/WBcNTUc0QXm2XXt6CVHUg2ysNQ9otwkTHId5eJ3NNsDQQhuTlpAsIRFy6mJHYJgKhZ7e1
BIPUGoYOUMFshiykCOxeAuX/VHycdHbfXitb+X0BuBl1+UhdlCG/O0Q5uAVJKs38QuPwVBpvYl5E
q+mu6g0hVOwcmtIYCfjHeqWKvfJNThz/gjMimrPxUfdcFkRxyxKa+TrwkuQ1NuSyR90qDsDW4Q0Y
5tL7um4GJ3YvWfuCn6c/zCgOABCIZlfRNSvtXKIMwjk36vgF4U9UOI/L9PitsxrhDyKTrQYW5rAP
n4bW6+3P9x/emuD+H2PgInErQOV4/vxJNXf3iHcnBSB3rnO2N3yvRQmgO0lSBF6Vpk4PUX5P9i8L
vZ3MU4z0QFqU9gTl99jkxmTV0PHZYeJAx68nfK4bECjYZeHlPSqNTRYVE1dgROkIiAryCyFjngV1
MinOKQcGDMkZto7WsNAaeal3Ela425EVwJ14ohwX5aISSTzAaw16lq4jIamTcVa/zmsHWWZRtyJs
5cLnZPfGS/S+I3n+gRe1r+mg1b3G28RLFIQd7IUUjq0IjWkkM7OwjGDomi2vR5ayo9LJzxHj7Jll
ftGRJdVsJSlPfWFmPEz2ozIe7k1LHR3WKmIiQolkOtbSoDEbqUOfd6dhP8HUDqpFCNsTMoQ1BBVR
dk28Rsy19DK15VWveJzAjoYdW0GYaVndD7HQABijJyaOmCjl1MUTQFLEQsze5vBXI1aBgkueF0mL
k5fL8L0ODghckjQBO3/a8KRTJ0VTmWRZ3bYz5baa38Ypg15u9FPBl3PkPs51tcgrV3oC4tZ7HD+e
p+ccu07iEfPVFIdeXL+slBdVA6hG0B2yqFEtbuod0GwwXuxebXkBa2tCjzZrPU0N/aDYd0TssThu
xRg2A6D9r5YOBWtAClbsn876/hUlnH4AravY9k4nWthSLxDI/nqN1Ha/soFigb23DFsXTq4DzoL+
JhEj2WyGeejY4DUMx2gSUHs3yV7TXiutl98ydCCA+VndN0ao2qcL52dJEY9YHAHZGj4ilrqspKL2
rDLo1njE3zT533ai2Jtm5iZu9W5jEmOe1PLNNXxek2HsBbBc11iagDib8KjPSfZywr5pTRRIM/gP
KrY6Q/GBot+ATjEyv+ZpaXU/UBR5NoBh/aKzGcqIAq5+0HXtg5Jlps/j19GUin4puC1aT5vJG6h4
y2IEwZq15kymmlvO7F6rYlo7aeO1lIGYOcINhD1Ovb1t3D6VSJEaRlADg42qzdxioDai5qifJT4c
MJA+1BRVXSL/vuRxKCik9C376CGmlsPrtb1NS0L4WQIVwcVkRoYxQFy7mZVi47xS7yqTXTlfWkyZ
xlX36UZLKDZ2tiKgOilUXzc40ufCq9xMsISn41o7aai6IgMsT/wDlNr2auJWWmNaHtoxsT4/Tj/p
wjcjObL2lTf8eDw90aDySt8EqSJCCiquEZw2Li1BjGxvSm70relfsn6+LdxUcYt+w8TsAeu8DiWb
05VzcZItnCIMi63WScODMHkaTMWsX8uTC0zvM/8q8iI59mMHRCN7WYEfXOPeKfp6Lu9qu2VBo5Ql
xCyJG/8kXfI0ZYpYnOp/ZNfo/5ObdudfUkNVbwPmZVDbea7GjQqNyKjtO1cnToXWbOmDSTHyOM29
Ph3phV1hPaseQ51oktDCJnnZYUcT5qgEaH15XHv1NTV9kjCUaqVUHJKy/TBXfAaD7RQ9UX5ddcel
rMCm/G5DaH9FS/pyvKryv2HHnVYASvjeK6iL6HFLTCYW1TY+qIBOXimwCSoExZQMCjAt0F7qLem/
n8Mqj7VcxWZBtRWPpprpaJDMQmsSu95ZotpfiEH+7PhpThp+r+LYtxGgQ5HAs6vWtBAdbhxT3oAv
+3+P0g1bqfq3wofakkIR+bMhV3oEWagw2/nt6jrB4YDyKInwvyBrlr6ZNws3aiPPVW5wvnfojMqT
D34mMMqdPt9Yck7Z0wXzDLJ4OKgQbkT5gGm2ofnGu3W6Ktp3lyfQ6WKAiEUTJqgWjnL6qUmsnRG4
R1m6/UmXbL8w0eDkul0ux2vnbIjYWyJZXRppzN9UKQ3KaX2BQhVDn67rTkdm4akFD9aXJIbsvmYt
jQWKJJtiVbDbU6ImDJowRcDu+sjYM/cUyQqdmGAJPUD60cDJibwPhdRO82Vzmn5rk/E1Cv8t6bNG
0IFJbgZfnWvaTiDLqUz73gcOTV2cV133EiZUHZ5xECSykayqH9a3ZdrzCIFnoQ041EQLY1p48I+W
/4Nq/nDofepjL6REEDbU4WJ9APHlRSU4U5liBq8CQQo7AGBxaPRPZKYWQe81+Qj9c7AMRvjJfvfJ
TMaRSfBOfDk8BO4jv319BpKHqzgu2hIjjN89IVcOKXYVuChW9RD+kzSt5DePD4PibWOgejh4KBgz
ZC5fP161mWOwd1FmdLh5v52mKOpfSbImwDDQFgNUA9A2lpq3Vr+JYFAzAQRNit2uJ+dCT7vwZKVK
jPwk38yI1DglnBMNoy4GlYoiJXNQH3Xv2QxENDE7CxEDy4QZvpKdaDKpRmECHoNRmGmy0iggLuIC
z4QmxIR9b0vVs7hoOP80WkUnzIFSWFMrhobKGxAtdxCrRHkTCNjzSMniF+NGlwcKR3QF9HyhOjCu
NKTj3i+58RT7Qnzd4CZV4BRq41C1c6TLTQ8TGSeOJvDFHLgNFTiqsdgXxNqVdMN/EY3xzRb0M7hF
jSEjJfD/ZJ0RiJqyzQJGEa6BrfvyQA0feko17CoGM/2khsIm3ZFB1UsfAhzhvVO4nlcZQAiXuxJv
UuRwnwSLsqdoPrInJXc9uJlT/N1xeD8Nwu5cNDsBHSENoJrG2Nq/f/6AOQBWsSnHnm6csyWzlf7Y
OeLRmL+12sAv12jl3Pi9OhXdJQ+9pj44e5l9vpdnYwz/z0lsjWGmzcVaqM13lWxGtm4y0oaQ068s
2jSLZTQGjpBzW0EnlQXJ1MDhDeovbPz+JRaRDLrR7EB4sbUsvBMVXeae0sKT1MQMqTtvPGZF2sHX
c5Q5FOnTLxxHBIN0OYPSZjRA7j/veBQH9LO6o8VEmFQR16W/PUSQ4RwSTTMnsGW3WIDkG49d6eKe
lyxXu5ZwYzE8jOgf7bn5NBHx5Qjf0RBnVTgqDGJvsPkgSv9RkwHijKatsOBwJze2RRenrecdXD8V
0F2jJzMeocFDwgKIwqsXIUnct+xDHnkB8W4HsLHElvezEaL7HGp8cGUYAILwuTOFvJzqNVCwRVYT
8KtsCDvoIhWc9DcBQw+i5gsEhD/dYGajnkGpaIqGi8MtSuO84v5geOBAzbRjnUHMLeFiduBB3s4b
UnYLwSzH1bu1psHmeS9urdci6O0eH85ilecpA8YgDaolrtQ7YQGqfeD7MFAX8Iu9Mas8zpP/6vwB
59tmxvTtSFYpZWWAbnJzlzP1mkQ2ZFS5a2FaPjMschWj4p6ehwvuGI+36+iciJ/64XxuWt6GXGbx
RTyq/FH6R1xsf6xcC7YfhMeSLKVYCpKV4rItc50TwBYEw6kkc4gKnbNoa4+EunSvB1K9+hddN7R8
/loGLULGuiChkMfuJzyr/N8KJ+vSGrTJtGQu7tIjuHdqMtI2ZQSP3RzqhQ1CwajJbZH8mEP3CafK
ahsLrG1H6c8OQ46fnCGxD9AVozXwqa0NukpPMRDKj+BBiuZy3FqpuQ5DxyIXdCaCbZPuEReTJRou
7trGJEpqVF2UWAGRvJyaGFbA1aQK9+9ILDm5zDzRGVk0Uxl7euXTyDNbmo+At9FCIlCiFAHCcoq4
b2uEGEGPgEDO5QJIaqqKP5EcZFEzw8yuPctVAaZHbpmRC4xKY85hguhLCdfGW35GpMbRYzuv0Db1
VvebNeRjbptN2Cg2J9D25mYJqLGQA57ieEQPxcdt3hxb+1IjkQAEoxc3Jw86qCDT5lnPkHSanXaD
C19Ekv6uihtFbzTv8r3wn0Cb6BBCyhUSRp7k8c7oLfZZZOQRsgMrrUyK3WiznqmxOHc7HOfuFNJU
CpGhlx+DhgDBNzTXdVOWYac+PnydOWjHuEzEvBnC6OPUQdfZ3GADRG6P3QpMpeeD2OCuVlpHcJwI
c1qRB9a4hHST6goOGNtt9ygTw59SgC62pFtQn5jTg/kmJxxAYzm0RgMiM559BAtg0DbzTAWTEwf6
2ViM8jwaPU2v5W5EZ4Bb7qJDQoZn0VDH8bGHIyxE6fznFn/JMeH6VohIFb/FydjUGXzXrr0f18LT
6ByqomqtVAbsEGvsd83DCv3wr+kWmMKqcbOOCgvzxM/R2+2IInx+Tv5dDe3lPxt50r4kZuWw8oMF
HGRSKXgqPkLr34PqRhr7uGBOIG13IAiKwpA+LkUKO2NPBw57FnzMslngLTwO6WHJwnhz7pdxZM6s
wtysexAxiBIbmZCKspNjQ8QWtVD+a1poQQ6jDBJ6IkBAxtQEcvdtzksZ9j8QQ5Z+UZUpeiQpNgI3
85sbnbs7hisV+Lzer0BaxdbKKgv8l+1K9QtNs1j8hBlvNQjUxc5cCj5piGkZnZLMrOYkGhYQ4Dzz
y2brep/edJ7rnTJUOtx1nB+EWd9Arr12s10SvsJQxPbdSjcakNHYz4f8qFE3mR9cEFj2psFym8RQ
Tcu4vKs5rgLEvq03H/Qn2K/SFF7Na1q8+iotCCZMuepMACRKDPPOKhVBkqIRKVAA/CfD07EmQLQM
yc90mR1v6z9rE86m5/VH/EOaVN2wbZZUAnVYfKweYVJGfj2VDKZlGm/QleOyHlwWXxSxPmuYh8c/
D3dmwNPoe6xgijdAeiBMDVVXXAuJjHcRL2i2DorcfuRvW42bASEeYdnFn3n6eXpquVCM5jrDeDmo
+XeBBcnEd10P5V3gEIwAyLylv38T0a7eAyNxGyafWkawW2ES73dP85m4NfWXjPuerPRiRduBxxIz
6j4f6OYfM1ipAJthGo7j8kOzeyfTKo1GwDW06MuWsz6bRkNzMA1PTt2jZ03m7ETpNicbK1cJ6crh
azcK+VhKEwm78UCTCA5pGRW07Pu6MYM+iKs6pMeHYhVzr9/c7zZIycktpuf5AMDRjY/zKJFsV6Nn
p5aCq8OAb4MqBBod7ev/tFxyexJYUIZBSnV1csVl/g7KNHNq4HD60Q0SYtLsMsvlsPV8+tZVzn1m
R1pw1rXlS1NVQP7Q/Iatte5s2f7IeZLQXB+pFcqupISjqgBi5D4RVXKVDE/jTW6IKzGv1DwnfQ5x
BoXII7Pcfs/SXIgTlJY3Kmc9bR5lWQ+SkMWdKjUQGv/oAv9tEAqNk905KMD9rguLx+TOGdzEur7v
xbdZhTSfkilvwK9Kx6e+HVUZd7hJmk6RPJnVudTUkPveJ7xLglU54yJoN7AUNgh8hVJshs81J1vv
C1QH54SYDIBI0hrH7ybvqOwwtMHmSTU1WpRaShCHSDs+SgtJwcrA/3fS30qx3nxxXDHDXSAVLnU5
JGMdWSDq4p7U7rKVmBudZLGVOf7DFfZgXq7+5VEOwNbPzvA1xGX+6XUaJIneafhZCF+gAP8rArU6
V6ZutuUUkgOmVEfrfCgeZCz2VXYHKOUHN3VB6WqALiWmjDjPlq/W+JHXpdtsdzUC6yDxrBaC4ebJ
sFA/7XHMMiJfzvsjfOzgF3qsYf1G2FSxLZTz89Y6gxBKa24Rx+j0nLkK/b21xkyEF+U61e+fAByU
qvhV4T7M7btHFo/SVXNl0hItk9C+XPEZAN7Tj3MG3NAqlzRTwfWkO6frFJFw291LlSL6jouRwk00
w47RXUBV4s33X6vw8SUZmYT8Kf5xSaNt1DnT5JyvvI95FiVXitJ1AiM9RZ2PZ2c1Yq9eYR3VeM6D
gjHPs1sX0Gweyo+ASITMa3A6RaFixkIdahcsnXJYkrz0IXo9HBwPjGE3XxkLTawS2ezECU9rPQI5
NegNA/zUdlNHa8Ac4GsJ/CkyKbRqXNhr304G4O8jwtzylUoadAkd3bUnf/D+vRMIMvwWFBPOv5Ci
uMh4YpoZNH7sz2lz1mz2kHfyz3MlfiIannp6iDxGXZ9on2JJnYancdtedpaK8ttt3hNFcZc/+nd4
bSOiwGO46gQw/90izemi7VaYx8pnEiM6hOwbOwxwJo9jka8p443TmIT96ij1/g5rrojK5H3UbD0S
sh/v4FZwub79Ssala/scGnSMIouE4bOuSybD03nY9lWuDqiXT2XMMkv40+DmgIy/EmboZm7YlFyG
Aiox+CFkBQgr3Jamug8m9b+S6NcC8PWDOsf+XwZ9aA8bWPidUw2/Rwsj69h1WB6T6HJRSQeFOyO6
aqYAnVCcELJQNqd/HOk/DMVV+msOGEf+fy3Mx2dvEI3LxxtI6ToxxlgLH22j0oLE/bS7vmVZm+WM
xMgyOE9db3JTKvyzHpqSpVQ3tmpWlslivN45BX2+Vz3OFK/NySHe0wvroNe99cpI3uLwYyir+Kej
SMh6c+1nYEeTlOxKP0EgX+QDND5fLbt7oNtgUS7vCp4NtBJHRd7nXZyBzqgxgtiEaasqBjWDwOYn
+gGpXmarS4DlcSQmrwv7mdJ9pc0M+tWR4pz9kvfxHw3s6nzz/Mgp4WiVNPPXh/sQKoH0mEpPJeMS
w8Q4I9d88ehGz/z1TpYwC7XsTJFUDqA5hTYULzHIvC6OxNlXOQgG69joQvugX/QZO0q9M8DDLaMP
qGK+tTxKqktr0opxlrNFqkkNApFUIYuyGLhK2iLTqrdhFSDFN5RE4dpcRQgoeyE2JyEWMdqo6qzs
2eFphS6kHNpnNx5qmP+e72ZoC4DA+y6s4gTMnpXxU+kAvVPlMI4SNMPrKGsSFYIue/rkQ4jQSPyD
CZYeVJmDZkhOItKtP+jY1xtha8rw2So8MNagaXEKhCObHgPVoj5vazU5UWoEde2+uu8VjmeSeKwI
+EGe8i8CxWVBlDA8dQblR0LfAMsoMv6THbRPJUCc5/0S2gi+lrn9bUqa5M/rAhZfI8tFGmZ2dzqD
78DxIF9P8fdg9HTMk+MlolNQHDRa4thuJr+7g8+PBGX4azOZ/SK16OxhdkyK2APIEOPntoRNl3/u
1rqpfTgdJtnzexVGtK3iTpR4KDO5HYS13uV3Cecb6VjOnqAlhpdQ+mKNzcTBDf9ws+J5KKPQtFVI
MMea6EVfPj9r+/dKng+oxI9FMRf2BRLelPZQL3kMlMfF6tMOWJ6XEaNQRMZq0VfD4B+O4HTCGhRZ
QhSIpuZ39ez978MI9veZEpvnSyARXRmsZwZ+k088IzPRhwifQsVnVLdIpjGJbMWoMJ2HDxgsC0Q9
vprUfH9/zr2tipIIAn3RPAh/LwdKXHWWTJRel0QZESrwxuaZbc2C+yZ/kXVX93Xbwz7/bJsiWj3K
vGaa62x70Rs5kpTw9dGa7M1wUA8Ig478lH13q62gG99pt0zfE8jz4JO2eVf87x+MY5kv7UshJQXa
+nAtpAkWfR8m3l9NinyiwXuaFdKPtmF39pK/8zQ4h8MF8+2Ol2ZYFBqAcBLblT5M5RRYQNulEkbK
lvZA0g1e1AK0nPctYhPLfhLYCs6Dtlx8iWZ3d+LzhDH9pXDTQGP+i+bCn86vr6dCnn7QGdk9Ogc0
7VK57gxx3oAlaSEgXQGo3oT4icoYdbjigU9NzTI5ioHD34HRaN7arWpnlov6sbybqKLf9KdMpHMw
VhSaus5ZgFdVPm9wzuEihMt5QP7o4/T4Y/u/WvvSW/jDxdKuPCaKXsKobJo0qdkIIFD7YFZR1lxu
NMsUczRjWJFFfl05sCRhB/rVUH7lKdF28BmMh8GOVVkHyEAY7CHHXWhCPbI9gDVh4zHZ3Ddw7FzU
iHnjqG8tWDIQBXSeYSttSmHywVFx8T1SoTIc21WB9t4DKt9kTgZD3r0CmyZ+b/Xq1U25+koMTeE2
hPjj3vo5L9Fox9CJb7TYlobFc55FTCXmKZHmIRv4aaSmZF9lOFNuCr4atr/5f3gaqGjOhpucImfj
S3+Oz95lJTHcs+158mAo48xKLF1Tc8gQBVm83XKFmBpSsRnF0D3Ao3SpP3nYMF2S7nQa9id3LAyW
rKUJB1DT42DRNfwzLJrxtkY1jy0FhpVkfmQGJdSER3/0zx2GCGBUue2V7++0YNm40CAaPDHITPDi
e/w+JictQjm6+SBAx2RIBopgJg0svGITOghasDEWgNDuhMUnVkK3wtpBQLwOGkXGSYzCpkblospI
pC8YpqajWrZnq23qEKerUbC0lhK69NKBc5p3RZvviOhBfZ6P+fIBsCDWlm0L0JVWG4LRqKlSe6/e
i4ownds54m24HZyVxXqeALNavMyhi1Pec7sV8dbOfsmQ0d3j6W6I6wtzHNjhOM1svYADvwGkBtyS
E6wA0S7xGuV+Cdm8/dtBmkci++RC/wzl0qPRDPsEhigNBmvUCICy65kh74mF8FNe8bKIL2U3Eokw
e2rVCItMuJancRugxEdTCsDDlo8V0ZQjk4ZIoxQRVAC9ewJ4D1I/M6Kp4JXcPZQnXvdYSk0HkueG
2RLigUnZD7HjY9aavOdMztwjPilAJqqwa1tz15Ui/kTfqbywZHupX8S1fH9bLGseKulGTrXer3tk
iOtP+lzEv9O8E6mBm3znSd+NqLasQpatbTCJbIVCXppWZIcDG0MbDtzgGCA4wtyztJwow+suyrFN
3AgESgL+9w2rj7gu2fcfCdhABNfWEpKgHOQ2BmftplN/brBKEnuwA9pNtZxWJPwpEojkYJEh82zC
FJMJ5ESHFnTDAnoMOJiaHzHb0MJvaUEtAWpno4GluKkXJHfVvU8eHm1tPpgexwbDk2Zf3t7yGOBL
4WlzupM/KF2jSCoViuWWKCJSdPP5AcAmSAwy8MQ2+a2LU5DrNV/nVvwdDLTUVwEQMY5k38LMmoS0
YK2pPL4hRICiIETop9MZ+IU72hWsVzI0tv15XTFbsZJV+LLlt5v7rQHp8MYOa1MXtwEcuHQRcbea
lzBuNyeTWanJF10wIFml8LN3iREGlIQpXIljxrbpyUPqjRFAIPPsyNeLqlIf7kou++igXlWLBMUJ
Q6FqtwmFRkiRBmtQQ1NT246YtJ5qFMDpDkpHEvcPp5eWYXfwtUBn/bBm98DW3AFOFgsCQzuz3SrB
zBvLdmgJ5bb6j8zd+MsSI0fLT+Tm+efrAlKwjXVR6OZ1rcJ6TtlycjFzi6v1ouT9UCwplzuOfdyu
KNaj9VJfuAN9WSDAP2PcuGL8mX28AtxzgL/dhuFssjgG/rTUey8diPiBlSIwxAa+ihaeulEeDsGt
J2AfYzsh2auJaNCzWljd66JUjEFIOpNfZt63CXvnVIyaXSAfssD+2xf5vIFL+lSMJvsqmSt6DJsF
m7OGFYk9FjDA0GQrWKqkHGAJmOgkLtlxYF3gq2x1Yq1GbEZdBb/4wiYOQklqi4AEDLiA0xSN01Xj
Bb+V9efQnEwtXJwyAg3/hdxaDsN/f7OutcQO1gt3xUIkos7LtC+KBBBN+h78kIjPB+dRIqi9sge7
tBWsemL3NAUDy/Vooiumq3Y2CJR+CwshjHuA3aaoPSs/f7yDsvyjcdMzLCaMSVMFSDJCVOxUzooL
YTqZadmDCQMwB5R7gwhFl2YdgB5CevprSx4Jm0FLZFJBGL5Sn37lsLF+YgnEimc9YQKwWkwF30mf
w2wc34a48R0MnyHdLS7t6FnBvdvqSvDD3WSOMaaLVbPhwrXtjAy9tj3v71CTyLnUr34PFIVUtCzC
8VnQqnXpiYAB++32Mgv/1No3gXJJ97t1UiZzWuny9xmKl3WLFfplDs4d0iZdfw66pXViZ+zZSs1Z
tk1Z3jYFBDOh4IOzKkHcSfWmZYIxdQMnkil5xkkv/9lGhM1UD4WGPEjQlJqvSZGgfNcc9+/8MT8B
SuDB/weimmTQhPtUjCTbbqLpusCBQsZ4gfpjRJpjw7SXp/8wuW8KpwsHhAGBcicyron9Bo2Evs2Q
MM5dsGbZEVMqtgX7d1zrvUi2p08rPQ3q6tMjZiKModiKWq6HtQzO/gK3UDvOlkVWZ0jJFMgDXF5B
qtHi+402ZYDPq2Dk87dx48bLOGiCrS7dNcmMiwjbkIQJgMzyK9IuF9XjpPiLNl5QAOL76C889ucp
Ftoy4mBgLIwqYISkEihdRa0j7+B3n7aws+d0HpEs8tOUXRCsdUpcMzGXpIepxkAemELiTQozh4p4
OLIvVwUI0lWIdsFTxjzsGZ64H8cj7s7ihP/9TRppTFPvT1eCRrA7RImRPBNWw9BgYYSaFxqD3kXc
F7Uim/va5cxjKxiqvs/iglGwfCD5mvSWhvXNA7Xq0nUCgdkk5TV/Bdf3ilS9ggat80REvNRiTCK8
pRqJw0y3kcc36bvtWukYGRnnbgRlYtcEO/QMwppL+nhdBV/7oc6VbzKntUS4h6ZTzzBnTpxMC3iQ
wQ5X4Dl3q0OaiNKEbVYL1bJsNULajDSDRCqfgY8qLjVHjHMrsoe1MmYAoObF+mhK8lEEr2Pp0NTb
PBEU6q+mEtPcQWPZhms3us9iRokvF4QkdtrN8fN7X4UjPqRDfNQu895IjhG6ll0nLjc6NKrTuAZ2
6GVvLPSO8LV7Kh6igYLABF01IG7CJPNK367g68KUnpJjU0OKN/jlD2ZTyd4aNFzz3omLFM9rFiqq
/hupfQBQLcKKTMPNpVJavrLPaaoRt2J4hQieqG/OU1CwFZvlG4uuECKqTQsxjemvPB/TBLD4D2sM
C2blEdZjN+a07ESvk0swk9qO2a4X8w1cWQFHWDbGa3Gpfe3bWQ1ED9oMOvqxXnERV7m/6jZULTDC
C1/p14dpHBEN11rB3hJWRrczIw3APeffgq6PGH/hR2ppny58NuxAvJ8ZMr6Vt6LROkMuYRhXrTfm
M1ZKNVKn5t8j75AGpUva5SaLaBcE8Ng2QTjhlzgHDQeEVrQQeKEKufXB8uQwVTAhHGgUqbVd2/2F
Z8TDanT2U07Q9VgeCf+fCoL6f9qHHS0Rw5y5KN0COGbg8hnW+ZWRo5qpnCE5TYnsg8VEFSoSlCMr
kiFhNTthspWGp/wwg5SCiR0iBRX/4Fm48d90cSYHHWwwk7JizmoFxIbEdQj36BjCnxjknJ+WZcU1
Wa6+H9ngo78IZaDgy0r+3dg9azEkgayQXsQeFwxpiqMmuCUJc4VMCGEDUEUj8jNTG43QD2YL2SoR
FBW2yHofvggxRZQeyPbMMMu1G5U+apsceqjnCXiM9n9HSWrCl8VcLMdZnbL5/TCEMGd+0vG279OL
1MF86fxwWMt7vADZYPK85nsqUIYj3fC3FLgIsDRpGaw7aWvVbtdHx3+xRDBKbBmcQidcUKES7IIg
FWc9mc0LZtGbjlbnPhfo8P/HQF6sg+YOIylHb5sWPBRMRm5tUXDOV15aH+kBd/eC58eq6RCfjDm9
HpfphGkZj7p2V7M5/5dxOy3D3mSNNGmA34HdQphyFTm59M+l2Qrl4AKIEH4UYuGuKgkKH7x2tavQ
0lyaZp+a/OvxBJ+tEzV1tyndGbCYZMPX+z4TRW1bsPgUXK2pZnKjjLssZePpXa7aOHOiUqI4Co/A
o7EfMIpjPyUFpkqHadkRPHJL/cfM/cCLmovV575llekvYnzDZQ9o0YXtBxWjohfpxT1yDAZb57Yr
SzEfAxpUkWwEAZT5AE496FqOj+ZM9My44CvFrYLcOrIuMGY49PbJHX7zOGJtt6Ze0Jnm8RxgTBIi
zsLTuepNuKWR0ZlQ+JCFRFCXmphWdqk1uSMwctxPNJ8iOSzbkJ/HozLUM8iqQn1AwOp90UwhqahJ
zNIYTZu0TxpZMcRefvf430/nf13NJO/Xh1EO+RCDoBFPJ1mpEhUqhzaAgHZ73ImHDXOwOpB0s7GS
qMfxYZZ/n/fSzUsQlsi9OuxEv/2T1CspSvLHtjlBb+GrKBizj7Bslv+MFcIRHDm5H1dTx0y+yRPG
Vv+npZS3SNjVBkXmj7mjK1f0to+1/9RXU6l0jSeZyS76Ye92unc2ZH0SSv3sHYa5xqKHQULWGr+s
hp+2onD8wkL+FOzbYNBPsphTncZDKBHW+O1swUCe1i+TXWKpo6InX/hFhJ4hxeQDtUIsMpLomB0H
j8KP9cpSH3Buy6G26rdDmUge1UROpbJKWEA0Z2DXF9gDq3X0IPKPwSVkcZlXXEU/qxJqhie4oaCP
1AWEWFbPdTf3d+QDB0YEZiC3+iw5e0NJKi6ew8kTcQk58oYQt6vYD/sVSuCR3M7ZHqQabWDqNWTP
PKaBJleB8d8VZH+pkA2x1S1o+EhsUDnpp1QiEKu8o4O0+WhhQNCMbO14XD990xTU6wxILACUonhY
yFUR4eQHt0U80dTD7sr3DLMw/Bbxz4kFKSrlx3GSajs0AjQRxQgM6NgXtVtCsvsfyYPCWtyGiLKv
ae8a+nT1awyr9N2JVFxQbtqsCEf7x90NvsERcG3P6aGtqMQEQs6e2B6nT7HgOE4lJ64HCNFqi6kP
hDhTkPLhRyG3lVB+L/hrbgBy+LWatPKdZqrVimOInCWbhLQqodoMzsMsceoutWzvetMLbAmpo7VA
C/5YU50XOT7bQw3w8PU3eXW1+v1iGLXO+d/QZxPEJ9EHIjxVtpdqBjkfQaLe9NxSJ05ca1MIumxp
S9ctja7xQij35HwfDCxJ3qdMJ129HVW5+d3vOw3zybsTpa+CvZ8KAbegSI2tSbmRF2Ok+uxuoytG
AobxjRNyxEEuVwTfGQZRasAug4FuaMqFdVe7GUwBmfeBYzzVtOYAIICTFsI680J33HWGEx5dRG95
ygEPgFZg3yBOK1ENwY5TXpNgmQ83LuWEi4MgtIp13zXod6vSzIkzioS7ZYNs+LwN7px02uI5dpYU
DZmnx4yCxj6lOWFCb6+tZ28oRDdXvEdM5b5Uouh5FtB0z7m6GMfAF/3VdQsd66Ie057uhOc/uZk3
1O50fnFrkGUpkVjGuSqXahpYr18L7bcMY524/W8RoVTw/Q+bTzVSNDhPXd9wS1QLpyOFxlFDoTc6
ttSIkMVh4fH2ooZBaVa+PkLjJhZ+8ZwlgMSExZiifNsn38NgmWaUdSV8Ah4ubQoVe/oPTFWQvlAL
3S+kh83hqAb9VgJKwm6MePJxX4cgQ+Vrjaxo1xPvouZXLgEYTk1lMZbOrVpAUqg628prqHRJ+RRJ
a3VElqT/BauQ5pNBQPEWnfSECqahqyXXG4sGxzswk373r31sbs223m2OyLwICJz3P+W3MW+9fcD/
IedCvnQcnQEYmGQAxGnw4iRQv3WvyGRgbTXZ702jMagO2JBR5CF0FUNnZvvV35S/RT/zOOiqmGmK
MXM5QYi101ixSPMITXXm/f/Cvk/3Czw7V+5erCFZ4Hec3ffaGD/30DTk3APVWw+pPx9Kf/8fLrtD
Nr9cWtPQv+eFB+IW+RKeE8eXUoZjBsH2iyr5kDK12BJsV/Gc2+VBCVJnibPycZ4o9XFg7FaicrYx
wECQj8FwDtJS/3mjKur4pDmPp0Rm5XZs+mi3xibFtJI8YKB24Q82Bpzf2vNLOrmuXdYcIbfZTMzf
mBAoAstpOEMiQD+L33lGmArzwDqzEWwkgKElXZia/VRrWoYGJg3DCokDDHRd96a6AFrN5nLEF1OU
YnA3lZ+I5AcW4ZYSOcDggDzGA9szFneVCjPhYVraA74JTsoLPmv09dTT6dC5xZHU0nFZj/hAW9HW
N/HRKPXp/IGG27+F2hflAt9QNL75KamFi3UmxvpCWWg+GDwxfOG1CjvbtRLHb6vMUeT6wMgjdk9o
oApl3q6JoxllcD077lisU0o8oCjhDpiPRDKa8mUEu3n6K7Dwn8QvApRjvKRIfaQWWcJK+M+9n5TU
Lm48R8MdbOppXdeIhMdezCcDNILJ3+p+c3QXYkeUAgABjxkrF2KiZXNGU4bC2+K91GJmFJg5Ot6m
7YkAduEjWLP4g/bsWA4dVNvVbE0l+UVh/hG7baytcWkShPoGoIEgCtR2UPlZxyarERvW0YOYoR5b
+utnfQ/jZEbKax02ujpLV4jUWvUE1PHTSXN3jFLz+MCIKviheOJ20C3Mw7UmklOCXs+f9w9p53se
cc9EvcHFWVxEBEnCuTtLIec/imOb+ctJssLeEk8vjvqmUlgCM7cD6+X85Q89gkHalJDb9mucWqpz
xgjsgfrPLfvdGy6z3gQZ3ZBFvGZJYZA8C3nUPLRGTY71h3Q1s54G1bDdUHuWeBnH08v+9Yfse0V/
V1o2qXoR6+d5IR/CyNX6RoBf21lRGLKogzLSkO3dYW24TpiIB8qYSce/4JQWxqgnz/mTezTL2hl2
zLC4vPHqojR5jhwXusJHnhSEPoETtCEtlTN7QVOswxkozc650afLQgrvv2f7SQYclLb2R8b7kb/h
yvH6Lh924xhHaYbwP6SsDKgGzotCuG0BuCaEyQ3fDhQ/A1b4teZJugqCM7RSvv3ns/bvbq+3O5xb
EOCdimxlF9yEwuvIx1IlfGAcRbcp7Gy7zmHvO7nNAJGCAyjO0kEpuZpd3IRlGci5owO8BIKz5UEx
9J4jpjOJ+tqh3rE3ykiLUkA4YbmU2EAHMc4gcCFKSj7r1MvOgnXhtoPezpLta5suov/v8bX57u3l
MB8oJK1qioS6xnLinJqJQIqSrTbJl4OxFANncChQg5YPJXXPzo5MvoJ2Vl6LsRNFj+MLJ9B7gq4Q
8Z/CaWxj0+Q64Fp1UjsgbA8CL9tu3jCIPWVse3F0XKMBp5YfwWkfN/pqH8AZsKE5gpgJrX5VMkSr
i3pUHKpQT7d/NhNJjvq3dp5973WdIIU5wsDkpD8+yvRPW1aKM/DR8FbaNaePyG4PJtgTZzgvibCT
K9AAiEIR2LJoTtzNeAywrKX5cjl5uTSnzZcNB4EBV7PQaN8NrUWWpViglf+gR3mYgoH3CDSSude2
NrpG0UxARfU76tkpSssx2KUO0vQRwUtT6RJpNdT6KCGrkbkQYEV0/YHFmHgRWudLBn0IszLY+oZR
4g+Zj+RF+JReUZ8bIjssz2I9FIBe5W5ENOIMig0Oj5qYH8GbHiVQKVi9Bcp2zUIbgny8yWjL1mrk
90BqHLl7rSCyHzV5fvotBr2Kw7uH3ejjn0vSt0/DKLjzv8JAyPOJynAMBB/WA3IAEIJ6EIc9O1Ly
pwUIDiC2yQ3ZQJAW7iFErwoJnbnIQaaRN8mw+NfQixNInftK5TDyNeECSTRR2aynWRacKAzx+czx
22lZqIgcNi7SoJL+/4fKzHT6bBZb9FHe1qS9gFBXhu/EHygB5/kD4iYNxn+iItcaRaEirsXsNLGa
mo0/TK86L7VxIcjxWxNyDgRJvYBkiWgOyFUqVPLAvOfPRyhSY+bWl4zPK1O9vBw/MUh0l5OL5CRx
gFArysZlPxMNWX4Nb0tuFCTwdIkwJ5vmw5PygtLT5YhFyHasvP0X3CbRzP5RnQmCPgugjpS2urb9
743idm80MgMi5GA3XGGRAxscxUGd9/gkquIlYTsA3QEMCo+EiFgkL1aUX/NI1jKDcs1kbgRuIUtE
000pP5NGuFYbR8nRaWuqn7GhrCtq2350gJMrLSyoGuUTQwNyr/jsVv2ru7WJS5YMbmGlbSdhvTNL
IATinPncqHZQ3uMRoaixZd0ey3nePNXVa+cMOR7sg5x9NM31RNEd7y/vTgM32CsaqMfpQOka9eKg
1eBQRxJlUbbk2jBXppekE9nyJqjQnjxzgiXw5hs+Gj8l6A51lz6iOxUe3Qpth75IOkHWFb+uBT7C
8tgnfbF5dyOYy14F48OoIac7cWGpFz+ztNPSmkfxQ0qhfYxR5phLyZcCNVij31GKQCjqpG70Bwjw
Y1uiEA112VPOBqII0N/M3zPJPf2RC8t4TBBUw1ChjPRzfzWfOlXptSXdHR1Vlc5rfwH778tk57Q4
uhxiVKJ4VmNwss1iIr0adkYbv6gDYJcClI/wiGiluNKjadwHJ7lerabWSm17uu9H/wWw2SDY/KTk
doe/C9+dHkFfckoIPoF+1i1fxZeZRcRELfk2NNx0rbNmzY8sz4NcXs3McCpyy0lUWI5wQJ3ObN3r
wBzoiEZyVIbe/eVXIrh7fppwONGWEI/LyXps87jpQ0HtUQohUIlOegnkabRE9ABXdi7KV088hbBa
BVQprwYoXLIbQnJG3u/jHaNO8+ciJhbIJxfU1Fa7Vpy9DFhsGcGKRPOOh48wLHQRts+WSUcb04sq
H8jxp+WeGW+9V3T/qVGfeVSoSuCj4fZQ2mvqzrds8TKt8hwYSNYQj3bY+ntfTArhEkdR9x3ZOJ0M
eUUIah9LSHDXhLDsqyN06E0C69y52EVN20WtNxTwpWDk1Kda/z4BNeLehyxPM0xA5e7+ZUW6JAME
rCz2RRUAuIdncZUtCalMBK7SClAgn+kYORGBvuo/MIXQGeL+xw+bMezBKwPXhiRIcG6IzJkrJtg/
YNnZGfZ0Lh3vdI4QN5G84oNz+xn6qLFFuiSfXre8WTPUzdmQk4t4LPSCiETu2vTlQp0/9eocWL5f
oNuw4jWhHEKLN+hdvAS7fyS83KWhuJst2qpGlrSi7C2OP4JxE3TWw3YqHOGsLlkaCguGPb1q2IQT
6fHO+bh0Ifp6t5nxGbdePHdkQ6nciWbAvmBKtSodtZpWOvFgMCAyL78KGm4LFXGJHveV0OV1g7Sa
7RY+AE2N5O1RDuM36uV59kK9u1J2g+G9aCtV55PLTK6mccxiBBzJ35qyrqElrrKNsOG9ykgbZoAA
ogWjCDKsQUZD6hApxWRSvQwE4T8R94+KWYsFqGyuIcTDAr6LNK4fwfu07D+i4esoWmDUfMiAR3Mb
99wbZilm7dh2SYmqtWW0DAr7rf2eF767/N6H87NHt1+hj/pRIEhYKZHo6oeavZwuhG0WFW76/co9
UA1n7/QABTqqSfdDtgaes2khdQuvvUl9XxBCvG73uK1rvQRPSb6ygbY2hYT1rOV5XG+xJzlT/BOo
Vp40OtxobmIxYiKq+j++BllHmsTTMSNOg0i9PU+3EDVpe/ZGzAW3q/TWZL8Ymy2mmjE+qkVLODVM
QoWI4Y4/rRsuFL+yxjgD3wLC1P55ZZ/rXBnWBFk+sOo4GhT8I7wBcE5kkod09EDrbjdoXE0OvZSh
WCKmkgQ33/92/YCfXbTzzFMCmtg9//DZ5eXVEXq4i6xl35BCccLSDa9hoqt2Vk8IA82WhNqLIU7D
jbDphDsqI3ps9fRBryI2H7i/CUK+Of5J/FuigwWx/1VVmvlBxs5jeWuze9nIpMV27Pv+k1Foanqm
a576mTzxa58xxuiqF8foNujOVSydxyo0q+tvDy3IW3BCOyZSRLcJTietJngeVVxeYSb+eau+Iox7
5xPKqGuFzOcC12uk+jAYX+8RJ3ctnI6J57txXscbqesNz07f3kIyDr2BIRXM7IJMnGKXCt3UGRTO
CwCflLZ1Baaan9rf1nMvVw+G1PdjLNCNXodTsRFksKwBrHD7ddJYdb4rP3AR3WG+6vQjzds2BeXl
x28RGp3SP6JaeZXGySZsWnh6DUTq9RL/bheaAyk7tIfc8z5E07YDNabaLWhFPj3X57MVt0J1YmXv
VnLrvooFYxJv5X7yMkJ+b0zzatnqCxBwaO7CltlloZ4UHmdJ2eKgy/17LqWRUw1GfZ8+Cp8mIh1w
NEsGafgb8akLUHcyfyIGyeQfbqlG/eEQUosa1p2HXzaw2L9rFck3FkKchFaM2eVHlXizzZQWm/qO
TA1UzqQJ+hWB69HVM7QBDbHaGa63hgzoPYigiKfyM2g1NC4tx4+NmLoZpFega4Ou4j9mtBScIegC
DQoRHrmyN2MWsg0I/x/6sTO4oVdV/I4uAr6sNPPG5Vz1rT03XuKrhsTmxuEOoLI+vD0JiMuTJVRS
4elKfDewq2/abffaXBZqoCMP+r982+H5xXa44IaryzjsF3Z5FegSECLngisWuBPe4xh9vUyKKRHk
MG//9Ax8CXEi5+WRNz9pTYPi04YqMBU4b4wRv55NDVCKHTz4lh7SEL90BHeH+AgEDHUt0Fp4dzGb
WlPCwI20C1eCwo2fCFfzYkoQp1WENfsXj62PeGPldaYvxMjCtfpLjEvVtkzmNh25NROxaFYWh3my
bTthCXcG+c7t4SEA1bo5iYeuKcW40AGJojMBhsC5zP3pJIi97Bvwrcj0JWj3RSMmxyCzHlpIeyZO
mb4QvJg3ocao6VGMzkBuN9ppX3h3BaPpckNt22mV0PVA63tR8hTQVV0baspQjXVwQu0whmpUDAWw
X4YLOyN14CKfCJ8aPdQ43T04VNMVl7LKy+dDiNPZ1HYfPEFBf7WLI6+AHzPT3G6lBcxR+n3hzxLl
k+kjQhTOQM/6SVh0egQpiSNW7BkLAiJZSe2FWSJuVG/weWLp/M97W1CK/48dHHiBZEOBOc0w8kll
lrSMPTMOsilR4MfsZuAluQkrY6dn7lYTKj5u4QYhdoKB7NJdwWrhUrYoilFEWHKbblC9I3PrytQV
9ExNltD3ICu3aFn36+bsRjvjBB/SChRQY8qxtQRd1FJ+miflkucvoXfq8G4uoL76oMeTsGPZJuh8
scwwSNXQc3WXw6aNZT6Sxep2sSvGCvk0rQck3qNgzFDigQAWlWpHsM63h1u5xR5U5NMAmFulDfKl
r2QILm57z9U6SvKlF+1idg16D/XeiUer9yDvsTFRHqUmEUEKDJs0aF4NMU8EsZsp2sLnASbQsO+p
pWQ6DHryxStutJZVCTjInjHp/yckMcW0VEeY/u6xXlln1TeXwILDV+cJZjLklX6HpjKXElIym6q9
e+nT5mBcgRvhqswO3UqFO5WL1WT58PCbo9z5K92YNxCRi7tL+UtONfB9/y8if7ZgnKZmM/1o4WVf
g2nvqbkZLpnJJJBCbgcMcE6vrAn6zd6wMKrU+4Pyyv8YMD7aYSzVYWNY7fBnwixeFEg2GiojAkqe
ZP8YFDGkn2SF8HYyUHCzdTDSK+2eUeqBCIKCMoOKFQG+YJUxTFSXGGiAd3BRuIdHaqPkhsAcy/24
i5x1mmmV/1qkkfQ+GsIYHn5BDlOys4EGAAAzW04FF0pk4mnC3lrXtEAZL5NX8fmagKg+fxV/bP13
TEz7ql8CSxlYmz1SKi5DXZtE5heLrY1a4qKqgYVJy1laXvx/sWHEKsgkDqRyp7mcCvZe2//rkrb2
HlTVyH0fP2B8xHjFKz0PrNcOr0Uw+1M2Y4BIpza0vD92cXW3S6Ii3pN/5zbbU7foZUF/WZhNF84S
XBt/9eYF1xQZ8c2Eh614bAG/P4WfxrIc/dScVmN526oWXi5TWYL0xcu8uy6vRpaLNjJZ5A8Ok5cJ
c44HNZf4SntQPWM4ECO635GNoMsHDUFAQP5/2qv2klg4vm6SiJPA+vhHbwNZSKC7BebqKt6qjtXK
NqAs0BUHLeakCu99KFrhvTqLAl0b1Q9EkyCc0IEZDZ+gqPy6cvIgRfwDnj541LOv9P9nBupuP/4o
yp1CQWiU2q4Iv1sMuZZVG3AntOuLWxnuApGGeZWwiVvCrIuA6fnIbrpg68JJePilHxgJOq+88Lt5
hfoUtiAGJ/1b+dd9X0Lcs0PvHtCDMN1wpySQNWYC2m+tMHeWWKX8JhSf4zAkiGJhYaMmP6iVL1gr
aYgru6RjjJWqofs6cz/yLy1vkX3lw+8DiDksTSy2OB1J7gmQSIo+IVJNUN4ERqGKuYm1VBhDC78I
2waLKWjmXRjN688Yc444fjNuFkLpThcAcsuPwkfKhuMKRQn8F4nkzR4MvpHeKBPGl0CdUCM8QBo2
WfjPfIiwGUNONQvfqehnX+wewky6rC95zHwsVZr1FXRY+a8MCj27XOWF7o1rXfBETV7jAVmLtOuN
jkkE17v2A6dfouoevSkyimWTLZzq/MEfymhyYtDJeLbIpKj89dD/uznHb09LV/wa0Wn7yV5WZyuQ
6Xdg8Yj6N99YrYnMeJ6qLxgsUlVz5nlST0u3fj7hgUhgoONnsIyxVJdoomA+PmcoOrpuQsGmLK5n
AwNGkaaljkQD67fpQB/TWB3I3E6abZjXhRwBb7JQURMdl4LDsGh4+1A+J18yEcR7Reg+9dmK70uD
tDMSlEFkT4+lF/wjiG2bPVbYgqcVm3gyZQKcdQWtW/q/WPTAALgsZeblca39KvX2KxnBFwPygAIo
40wF0PYq59sK46qMRSuEArgKTQ/Q+tz2oosuslGR+2MIXEeE4ejbl6ru/CuvaIuVHKCzTd/WAS/0
aTcbGgDKCqSswVnVtwDOXhsfit7XzahPOX1HEmfkTlG4lgaXwUexsGoqWR8uhfd6riactDGVG/5B
ikuxJIVeBNfdFhpmP/P2id3loV1z0S3JlSt8VpxRT/dFlZahgsDKFngn6htU6qUk5xrXZfbh6P2z
Xwug2+ONYLX0mShAj1J4ukcmeHoPEVr19FrLvlSl8904HoOsZkzbrt9wLdJkBaYdxpNAkqyoS1F7
8+qW2BSbCDpZhNWNga3Fqt8H82Cnj5zaFhl83FkhjiwJPm6kwInoqL8laAgyNFVDycclWtuLKKrz
OgaNSz8TurrIgVegxJQ1dVAf5Ld3n3XGPLyMjiYGpIoKxNt33GdXy+R4FyOQCxVz31K52nSv8xZ2
ORqhobI9DNmR4KnN0kdkbeCus2qE995fHTRHj0Y4mWpagCXdtLup1gFDq9dMg0pMGmrLtIGNdw94
yAG9d1JH2brksd4eAvOGBrsVmxFAk5cbVcmOLy8ii+50iSrKntTm9Xwt8qhyb0QZz0KOmTqfxw/I
gwejwDNtM0xNhZt7ztTzExZ12gs5rEF+egJbZG1e57zLHjLrFfKzK5D8h9Psoji4afaqm90hFQlX
csQpI89Vl8u/3957aFIaORHMo8RMENF0BIM2yt88SYxyeYJTTENq9CRnSaHAidr4vbttlYGyvH6n
2srzfIp3G3L3eCF92MKY8tMdacFXKOyXMRlGFrD/IIchvCK/voRIJeWAXy94Sceozx2JChXA9ZsT
RlajhS4NJtt5Fb2Xi+sh/UzQtUnpKcsXx1HhyTqT1NV8Hq67+wHmLw+Eqnx6AcGuR9noQJ+qKJpm
9nSk08aysjMeC96YaChTNKuJPnEIdB2KvNAh1JENMwt59GTl5Vv8T5vJO12qlwu+dUTUvrtTqinR
BqXcXQtjVTxmWKTVv5ZkcRdR4QTUAXzC8zj2O4Ad6h8QmExB0xUNXe3Lj1kAypBKIKCyw9icW5Gi
IjX7cpFgzkfTdcdSZW/M5SVUHLHFpyoXvjbcuzVHxHauUNDBj1DFgnvYlfBZec+QoSxbPJqbi//0
BcUX2zaKxb5udS5gMhT49JAbgpY7ZSobUPX38cytPZtR3aUptKCJ5LtW0maCU/sroBMGjEdBa0k7
WB42wF+UmLMkKjiKyPpS3Hy8D1fNXR1hzrEch3B9lPSOqotHh2VVjysZpUGoPtvYQHRseBQyobCY
roCBVyCNogakGCmtt8SC4LBhklqjqXFVCZlOhVdwwxJ5ZXtef7nVXHHRRSQMsa6KG+7Zn/J/h8ug
PJeWMOw7DWDZ/Yunph+IDc/yy0bHb8r2LR3LdCMwxYRutiIMEXfVwGU0ZjLKqoGWMDlWwfxgvw8L
Uslh6M5kqH6sSv6xKf2HWzI3lAIrcUNMzGUdhnGX9qBB3HCsSf/eTbcslPRvlq0fHNtddARns1xX
p1ABg3L/dqcZvxJf4Phq2lUSZGb6HXpj3voQ9nlgA35SMPh8RN20W8LYX0Q9kkyAACLPxEVYTdA1
D8/MH1dbGFed/O2z4kfcMZKtE0Ngpxg23ar8//12rvKj28F5XYQxg4taqxxoTozOVpciweMzsSz0
8Ek2VEdk2wBzTZhESxxTZZ962kr/91eBB5VmdQ7NCJECrklg6gCV2T05qQnuV1RBGnZ0h725m9S2
uP1an/niJ5oZg81DkfL76JFWSAg+U1sDrmRBDu5MoqrhTrhxFF10+DYLbfF7G0BfEirwOOpooiFh
vSy+5MILZMB6t0F3Sj0noTMS8yksWfU1lUkqFOVa31tnCsNlHTuuJ5NU5KZv4W/hGerdEgA+Y5oM
1UYDmcWRyo2Qj+VGO96eNw9DsG7ohZrk/mTVhEqwTtQEI7FvVeIsqHXRcplj2gBvqek6uUkh9xUZ
suwSWeWJWUS4Pyu4wSe6n/trciR/XmqLQhAjp2hVMheoaWo199dNQVUT0SgrhEYpqubiYfaKL1Wu
wg08Gt8lsjw3BIxMZdcd6fmezq6AfrKdfTn3fKFHKjky1eHgnj2CWnt2gmUjqRqLMsifMss9c78W
XWgJogFdcWXeuX2900JWgqhjGBn/XjaaX/NYRigmxkuOvVboKe+c+5z67z8umLKK4GWuiVKcROTB
iaS2II9LZ1OftGURDVW1wbA3EZoV2T6hOIAH8EBcdQfG0Ni5EVLJQQBqflffAjmML9P0Gf145zSj
vEp0efuP+zIB2/HJeyGnpwP7bUOcEDWsj184E14AwYTHc5b76aCjwtmhcNYtC2RbBuSLm50bApF9
dNiXnjNurgxkmzcMsM1qDueEXGwtcipTLz3KAsY7s5Tu+xTHMoY27Q6PGzrQmHtfbqqyDFP614NR
sicg2nrvXn/G4XQ6dr2Q7nU13XHUyxmHL/v+4vBMoRDLo5BmlCe7G2EOMi2oI+gUTswVLwQr8ua7
jAKoYBvKZDu4dB3GCbCrTUuzjNibg4/0ga7BjeihSGyrDu9mG0QThhzHIE0fGdfu7iByJXZkrRXC
/7dIS0nm3lFLKXizuK9RwK8edJA7yAaDD1VPRWwSq4ltaLcUw0J18Y+rmG+Jghef2XN5UL8f9Pes
ooPlzK5utxoklfMCn6iO3SuuHINv6pvlNctU77w2h0+1k+VCvCPlwG0Wyc7BCBxkGOt2ZgedQpZG
iZE5WvuIFIUg3Bg1ulvMyKkzjj8HUEaiaPaFFLdQdr7tXsT9+vyJEdhfi0lYggBni0sBjXzEYSbH
is3MsrTMqqHMEj6mBwEO7dOAZiZ+Aw/4tLkE2JZ9nLNBUxOXza0YM3Wl7an6h9g40Nd3UbXsKpvd
SbTrIFitXkO0J/9fDsbsuuKQ+P/HgyWA2Z5009jLPzZPRFDCZnm0x7/XHX9tcC6atZFnHu5S39+0
bzgwIwM28PLJFlLzL3J3WnrIg/tLzgtklHrn696+WoXK6AFpTbfrhJTVWr0DcPFn80FKEyIqkZ9W
+xgg3Av0yESdIvSekCvtAMEcYwVCMkoA85iBx6iu9tj3QACZJEwooafS/qyylhgdLnOqRL/E7Jkg
3Maw1CXYlddIsKM25PRTGuKao4oDjiXZP2MYS8aq6UNfq2xG8JafYrl7rjzgJoLMF0xxAc1rgtU3
sttljnRopUNsth+oHTBuIuyr7vw7+PNB6MRdFJz3EKpwLfYAmX2tNJVU00nQLemeNGpS+Mf9zlr+
n3iBX6sAEZMjbb1xI6QE3x586wJ0mJ/Sb/AELD7v9EY4KfC/MG+ptjyQ96v4H3oBga6T/pGkgQIK
KD8kTG0pun8GP6rbRApNZ4McNT7hkx2ZryLWbj2w8iW+dPNcW09banRYkQMll49G3Wapsq2X9zd4
5LnYUFDTbmbHsk2qmSzWKUnnnLogleqF1zi3KSD7G/zeBEkN0uEfedidIn0xbomG7sysvAyAbVZi
i00bUDNauPKEHD90BNianfgSOEd0J7XmvBd3yv0jX3l8GY4phqqFxFMbN4z+JNF9lDlriCMPmYvJ
WkrU+BHGnr8wuszhu5h9moqEa3hMSRg3h2KRenJnU5crRZInqr1JOqAjJp3d9C/mOV2CJYBkBD0X
U6cjfhb06GPAuwMQFtZiAq9qYdrR7pKbQ/7xDYrx4YcoNCIlUj2GAhzjl7QDPxoews+42UH026En
7Ob7/m9QigVFsf3OH3RQre9NdTEGQ0cGWt0nKBZndipfv3Su0rb0Jtpaf6UmSP6ZTD6ucs7xz9Ux
V3V2qgTp2iRswA6uqxebQF9kewiEOU88spiaY+nZcPIE9NqpmizyRHPPFIPUt0wnaAX9ut0DCKm6
KGc+5riWry8iW19AtIPCGQaCxgPc0X336mP0MJUXNUZRyh843wIOaHn+qNtnIBIqJFepFrIaB3yU
vbEwjaEPxDBxOojRO7A4aiKsxfpyYDp9CInOkqe3KVB9PNIgtx3leklDm+TgJdA7yOILJEyKTrHI
SJu2rvEZymQNSWjuI0QN/XETCj8EtuVcGwWV5vX+2P02L0ULlsAeKEK7w3MjI3shIkK5v9T1kXfn
75CTEQT+jzLQC5a64rzk7RfAci4fiehjeAsMd9QU+M/Jfn9XnlardCkERwKNSAps8yGD/OvKUxoo
trE6F8yzblk0oTOmqD93HmgTr38crzPVXW/Q57wMrrim0LVfdNGEJfQzhKcXtE0bpiX4HVi6SWNm
GZi22BzK9BFORYx6QwvO+v4DsoIcj7R995fCriz1/UYZkdamRVjp+WrTLqCl3IyHhgM//J5LoLzZ
yt63K03bv59FdTn5C5e3DBzjqz36XLXN6oX8FbvhDp9OjT3/QwTUfVoS8F3t49EcwT+ekSVmk/Eh
eogPviH+NiN0Ui4swx/lwcJP6WvH0/Ybzm04Y7mQWdsBhUMLKqqYjp+V/IvHW8MjUN0XQNaUeILw
RVnyEzjZkv0FPcNLaGd/LDdaXJ+BgPhx9EsgafHyeSZN1raNbQK/50d5EECFwF/33BWsfKdaOs5A
0UjseGY/I4IMC4Vm9Q6E3FufrlXwFIoN5ecn/Ib1MpH8pYnawjeeJ6GSJk7IizGWU1FflGyFmBQn
QUtYhg8o4ZtgccIAmDRATLadGSsT9/eK9kntCCov1H6TN9/RwUiJyhn3wllk76LkA36SElZH4iar
B8uC4XBrYCfIiTNuvZXsFrvk3HeQHgtHBA+WlrSurTyyjxUsMpXVNKKXrADdfDeybSpZuHmTObxB
p40h5fNHJQ4IPs3J+WWHksrdAqAfU7ox6bUh/THfq02FFGKFIquC7SdbWrQXASjJl8iu9kSZ0bBA
3D63l9D1wq3VMhSzzkIf4Xczg+XtOVGTlYN+3PEC2Db/1AZR4Q3hiaimEhD16E/qvj4BHsqy93uE
9QqpXQq/fa+8B+lpl8QSY8VvaJoJ/ojG9bp5k5h6iohe/KvSIAx4SHn8lw3lKK/S6WbDDXd154np
BgPiFIkFaPHGdNsF0Qnn/2ARX1vJv5HCP/Bs/LiEvWCxVawuJJS82uQLSSOUfmSDCXoFNrZWR7kt
DP8zJEFsWg9xAWz7Wn08Lp7o1g/oUMh387zJqpHV/Q5vs0q/a3wjhgB9kUSypR24qMFlweMmNSlB
VfxGZFdGL4bAd5MNGbLvXP3ZrUH6PTnQvAlPO71JQw4fDhv7lSwz4HBCEeIYL47u9eIhS3VPMf44
TPwJsAcSzAXIVV+CeQ269+s/WUtM/RgJaAvvxl2BhijrCF+USAG8rQlwK3Msw3LucpBXRgDONMg2
8lAuuiqja+noGQcoJ6F2/LgU6Tzm0yqFI3Vu/p9yM37ctoPpal9sRuGgP+rWxEG8N3a0XOVeZlCQ
QyB1SR48HxprkI7T+HxGt3wbFjLmnFZVuCV141lcN0Lrf+lg8e15o0UeqD2tkNbSQa/PTjD+m8Y/
4LG+yWQ9easHRiv3UilDLEjb5+ZNaufQbz4Kz2TJLlW1RUkqcbzvoSkwVKYrqN283V7LhEjaT86p
XaGCIG183HghHIuEkZhxY/p/De6o3bV0tH1P9G63s0Ku2NkObEqkx4bL+DJwMY2L8o2czNOWa5cD
ntidpAEQGzQtSJyf8PpcLz9AQawt18MpzPDP9yaJzE+3nv4T+e+JH5nXTE9kQTlCvFoqeNW3ppN/
oU9CmpemBGfCxIZprbNKKRh/7EPGAZrd2vEJ1yzw58TJd+d3sohO28mPVKawWV90Tl19+gI92sVb
N5z0M8gRdwXHvot+E0PgTwnBNAZL9+75x6PeNb7UnKUYij/uvGvBJPodGqByzJ3bmVj8oGEeK9Ds
2V3IBYhXy1yjCvpOMMXCEM5tKMW9vk/ELzfPTl1OFlp2eILFWozV2eJMc4Jw3FhHTjpplzrOdxbX
NzBeDT7LrV/fGWtKdLoOfVhwrcyvZqJMMEdiUDMlm3vmxjIRKnft0fq9n9SP78UaA5rueGmIVPnV
AsXEoLUquVsSkkEt/XGijBlKBVjq9w746IVkK9Xtx95k4UQ/f4ZhkxtS+4ASSfTJ3udrVHgg0KCx
r6eA5LoZ323yUTf/Hd7Vi8MZc6TGgU5khwmslAa1tAEV6SYo7G2b7hcAnTX7lGL0JIfzfoJhQXs+
c4HPDs0XhfQQqwV70ZOCl0voHYTu8xM/nX1nsLO3wpp8rTmsi0a0xwTcM4kcdbpenM2/CWn0NDS+
bqV+dzZQ0z8N1/5eUun2dWLtKJzoVLPL8PAYj3bLwBW670NVM5Z2TFNAwpn7TYHITvZqg7iDfUwG
oFOUFOfG22GBHoDyBy4rcuFjVqf0KUD2lxwuJUhlrmGHsGWDBwBofFKPW8Pvn1tmJ1ZYSaDIk3LC
wwANFJYgKvHZgNUKuAGvNirVZQJ0vAIWjKhao5/VF8hg5xAR7dRbxKdvkoiuzOEjoSPyYrC2TSbi
4Pyc3R7863Zul+7nP+jc8KmJza8gcDjNZVZjDcZ37ckPhkXzYrHG2FnbI+boTIanGyF82P/CIWjj
MCfeXRMQlBK95MVVCUhfjQUK/1vRirBNXAAyoa0BWGSPERKtP8FQeL3O24eId8Wh0RTcTn5oMBme
s9XVWzRbPahwnQnmwmgfpytYvcJFmYb73GyDBIqAq6sjybUvF538+t6c1RZjunIttBx/X/rMm+L7
H6/hz8oOZqwPAH2Qq6eB4Uaa/xmLexzS7da4fe8zVkVmvALTXS8P/sv/Lid/klNBVQoYYRepfRUu
oM/eLAlGSzirXpouinpOCCkmATdoz0JivKdXfDz2LPpZZiafuZ9lZjE3s2xDU+0sBxLgVVcufkyx
XL9nG59CWIZV1qBlHqIWPQDg1sJ5oGHkVgumhmUuFxRhT9x8NDezdrmjiUp8bsC6Hk6LCQ91jSdj
kxrvsEu8zuv9oYT7Nyl4MnMWkjEotyrsp8MPABJ4lqT1QtovgyTvVjajM8zTKhLlZnTjwqe26drI
eU8d7wFD9mPQyiwWe+gXbNzLTipTVwFBlnnk4P2F4hxyIB/LSMsg2aTomnrBG481SGM94s+wTixE
5ijxKjj9Tqu1cO9hl42z+6nX6wIUVPGzvSJUG21hng0YPBiOOwSwWP2iQ1iGSRMh/j0/2d+54Ngo
O6pArp83vx0UArYS4DDP/mlPYQ3Ei4dffsJ3Q5Hwd47m2eNbew4YjVhoCIQ0oRtU9/0MtlutgUMn
usQAyHji8OVIt1Cemx1yDaBWowka6UUzRXHRhmKRGlBLJfpvtr+VoVVId6r2RAm5aaAgStpevZMl
hrfJuYFbAqMHNKJNAo/N2pNu1F5HLoeMZa7RD6+GWsO3k2I+FnK7c+WcmGjrhWTsGRZhZ+xCnnvP
WwuyAjPS95UJU9XOucZp9vK/pRrsUS3o8JaYMlDeSvo3oXZPw5SvLYVDlfiTA40fahuXbMdibTru
GuIB6ALRvkTbiZ9iOf1xnUkDhhZqJ09UhHqQnSrIPGU1EJKO/ZzLdv7Ycs+9NRNuUt/JkA5jAYC7
IPQidE+GRN16z7zC3edXw8D4LW/kEdiBJlWb/eWUodPP7cGJgpbciwRVBeC/WVPjINJCpnuZpa5E
B46KPrx7523LuKsht9QkjXLiPkuBheQDMEx729rdggsvgQW6cpWgZ69oNpDRlltnb/DHA/yxKQEo
wY6qzgfE5DwNZc6B+wfHgK9qWr5F1RXLQb/uy3q98RNFTuQvUM09YAct8H41NGuX6dhc3jdViZGm
lIWIMLJ/wAGGtye2Q2GjRQGz4LWZhX26S9eeWH2KChSfCjahqe60lgTq9a8jBbF6O1ymXn7VDOAt
sQQ1xiL4GYtKIg/9mMbiXZxZis4Q2yg7Jchpu4UZDPE/yxvb6VR4o2wnO9/p4FUP204YBbo0qDNv
AEnqbSbbRUCiWFAKTLapOCSlLHR3CyN/0FMDeIcxtyiRGrLEH8/SkEnduYXKRq5kH7ZIcbR1U7O7
8qXiOZqGOx+j9uwYCEwu5Lvgj1zRRSyZQ9vzmDX3eXkOcnJxIQudoOqXySDdbg6NtaTxPZIjwURk
votooiNtnlTveAZiicpOe+tfrIm4SERQUrRwqdRDJu8u/cvQGvMyHcn2S9ImSXrHPmSw4Q7/4BTj
/OZzTaOE9xN7crWHNxRxWsrNlhZ8hJd64d+JR8YdQjnJmvRolXKWWdFnYHcO4PKmJwPlqT3qSr2u
2eZKBhbtBeSvRnOakaQ+9guSBAU2Xp6wDCB4o0PySzHnGXbvzPeVxI/OFvp7vUKOiyhd3ZbYOnXN
vbSmzBUDKJgM5w+xwB1kua5apiH9k5XsfqGARJAF3xGdcliU2RazrAtgvhNKYKrRBllvzXaLMoSZ
QZTvGd3gnwgP8uOY5MWjsO+wneZtUGlSFKbUdE2Y1gppqr7ckOy173apKOqJD+VgYZjXYlw5gU6c
fJkRl6H+TKfqSQ+IfqIdc1uclOm/WC3IgX2yFeOepTSmUe2+gaM55hIWpy0OZi/gMfsJ5yIhfx4M
Yu0fBPSalokRsr2Y3uw/y1SQp8I2+GK9rRpzgiTAmmxFFs5wD2k5HsitwewVgKkpS87kNJSr3Zap
fJY1FjF/G+QM5/OtsXTE5wrEexbqg2aMCy5SEVnVBKE84+7YInxxfOvQek5ILl9zwJvW/NCHbRpX
K3lvqI5xRceZ6E2ogc6yy9IlV+NZ574/pG00US3W6Xtzx1T7G3gYzHKcTq8qN4LU1DzcZ9RoFQER
RnPAU5j2FCyP74eohwCCSBJNPd8S73VOSM/+zEzgX+Niixs2apWAWY+SWvafZB9PQJOOVtBsnoJ6
1xUxZBnx8zjQGXqlvrkuVSRWZns75DWz/YyXVSh4UDF9ftu0wLnFQZl2kXQwVFLCAEHugWvjr0mH
67ujgZnsTEr4BNEC5HUeb3AmUGWbb0OtWyP2/lue4W9ILB7vs26KeICuRWZ1UuOaXkKRjj8Yn24e
FVmk/346sfUY4KFIYQszZQNEoYLvPB1ynly5vbeR/WnFTEVQ7W4DSqS/eIOnl/iiuYNaA9TlPsve
JCpYcj6MO8vhYFZaK6zeXOz1fgNpSohypxj8SUUxctH1024EQzRxBbwj9IexRYPjDXSaj8hVoYeE
efK4spsjFUSw6z0z/OufHBN1hK/HAwochYctYlx9Cju72NfB59U4860f75wasa0DSedgJR23aC0t
ocCcXALklIcNlcUX27tesdhaTLvwgjgZ5v1DYASoCxfauAaLjvIwZuULVSgCYTqcTTwcwJ0DPI9A
+3gBnfzgsUodbQm1bMttzN2tzqPHlOIIobYxMhRfFCUS+bPJ5hH3EE0k/xV6j43s0x5FRvxKXnH9
P7LaBjDXFtgsnM6/6IV0G0FlsSuGQWQob/XtRb3P0bPa+zH7YctZyDIPYqLl/VPy7SrYU1poDh5M
QdEeu9Atevt2DA4ACkXrj2Z/dmK0MquxvT9YX8A2Q/u9yFuSNU+7DqETfEHsE1tVWFzg2SgGv8n7
0FVzz94TONwmNH5kjH+j8yUPZS8lBT6eNitUYPiRhf0E/nDHS4sbOwzXiWhNKzwa4L0490oyByMW
xRsQiEVptefK1FQMSA8SXmApSOYize7YbUNKYIdnZReDqHF4i+EEN3zEQcFv3P200asitOsio5y/
Z9it+N8moUm9M76DF041fNrGigJfmFdjQqqbWcu3QvX0muSVXtiPEl/oY4sZwlIRyaKoL8scwUkb
a3Na9yxHtVM4a8ATSeVpYEuNoKi1PUS2SRaZ4XCHlFVzuiZ6YxFWUwfjG52WUN+034k2gBxfi2rP
30npM3aJHlNqC3sOpG1gJC0xTFZ4gTDKHG70HbkDLMDEmtnOunVLKl6agzGRfP60bMPtkxcJFiea
Nkbslw+e0fiF5FL/YO/6k5nOrlfvAcYGL3nVBoR1w7JNcLfCWDH3/4uRMrlwqZeQkt8I3/R+KHnt
AVCdV3bPa6JVz2LLdQLzssrExIOVm3+9DtuWSAbusG9nkZhccMyRmMqxABv6ZuGpaxM0ylsiBjLj
dBHc42PLbTO8GtxJvJLchs0/TncK7MPXeiaj3BciNr5hC1nALhi/bJoDaRt1ej/ZMaza5Zsmq0/g
WcEJwxCCXmLLcf5DDlnuhHPUE4m2XGF5S4JsNmdRT7DFRmmEPDOQEkl62xeazy0c1NxpH1ATBa1b
qPhMoROAYa2PqyaTAgGOxdquvncuPPs5B4iZ5HLrc1T8MahFRu3SY1SgrvO5jzjbt/gYv0gzOJ9h
BOy4Z5aXpsV/UGpdT5r6CmuAdE7oAWepkJsJpupFy7OzjEqscwbcLYrO3qkXX2wwXjit60rxx8rY
Wh4U2iF87xGqFoi0Yuhp9HNKj4cBO2nA6TIdBAEAF4bj45OneHSCdMUQyV8MDjE4WWH3h7JSo3mg
X/ACaWl+9xMmFrECoaFAZPAdbBtZ7PTAUQQPQ7QQqUYZOpqP7HPB3Ay1c8HjQYxGCm/c12Ovkf59
6yRXIVMlHvk43I4GFkGtYeod3XK94M7xqzBkAbCdcBKmjMFmw69dYOtR9S/xegUp9HicjuEoyM24
7aN5KA9yPSwu44RekjjSN8lfjTRQXeC4NmUyNk1wmkMGXd15f3Wt5oUo63R2quqpezzUfBIuconj
nhtmP5P6tjPi4CjI2JOHFA63aVocX2tNqdERKa2ZV02kPsVIT6e4pcjjKUDHjKzXcH09WGTiDRgc
j7eyIibhVDZwesJe54DWlZTSZQKehVe8jJHrbozRqQDKuC5AjPAT30rptgqD3W9N3hhYuUQSlfxY
SXaXU1K/uw+Mor1nwQPVBsSx/iiSPQvFvLPJzf3kZGhHN0BIZuDebJ2JwBZCS3ZNkE6PjlQdw70G
M4zUYw9QrFMuhEcXbaOAO5auWM5a6jeMrwx6616ND2zoJIyvJhQ6azaYHQjt2vPnIVeEjz7u6w5B
jJ+AqNx97irml56ShogWQWtzw5ohcZgJu4rhn1VhC3HqJPtcA8zTs/nKEzg6lNKJMMuyKIxuCepG
H4X3FAik4Q2JwLX1QOWwztbYkCGKRz+c9AyZ5eRi8JU3dcxAgyMOooY7cke5u9jqoA1Kz9539BXY
KAYTNFDV0pUGzQgXnIr9O+dNJ93SDufTO3bt6ToY0glxRSkkMSR7Rn+qnwNmjtOzo2Z1SRxAIHXz
gHRzUecxJ/uQerDxZOoUO8sZu9WOlAKxMDV3uIFo5Bcwwfb/ITOl0rel7I/jADNMLzEVnrdQ1WOR
X+s6fsfOtjtJT/LJh+16l/wrXTS/Rbw6jZTXKvEh55YIoegIy8l0scSoJ5+WhZlocZPQjD9oDQ1c
U4HXGjvrIAmPLVacdZHI/hf2XUsIZLFLzNhsMhANZ1aAtkW0qzMS6ZPYmkFvsjH8nrWakN4iF5WV
TDrQ0arUgr7PHjgwLiXWbeaZQx5RCEkxtAnyhco9iBSzq2iHq3Z86EYKJ+qG95uwZaIFGhWDnDdM
1XlYVprLdYYJjpZNUErZH2McCJ50yygF3M/U77rj9PjL2seTIjzoXdqD7vfWjj2KkoGCExFCGCdn
0Qr967YTfGBwbe0UDD9HriCGljEIFJGbtNdx4aCfzOmFCqiK1D2lFXBz6nUqL7ROagadjhsWHYU9
SxHoMrwfOmhYHmwTu5SylHDkDYjMjHGudJnFxUpkcvxXFvGBjhg9WeqGTKTWLIMBxZTgEw5D8itS
zNijrMrP27/lbl/zaEFlIbhzlWT3UFssTqLtCkm+36BsXYW3o1sLjhE9dk+fliB1UXvaW48ma4jt
M4Q1CJ+eqSXUAZ8bSVskVrYaP+oq2RTqn3KmLIQyoHM0y6tRo06I1FkfJywHHiP59Q7bwFo+dpUM
FEW1GV0uzEPLeHWa8IIstKbR6m8kD2iPdI8P5wt4U7fCV1bvHjofPvEqpVtRd87UbT4cnWwEMqR0
JzxPNV+ZlHqY1eAciUrsjOjiI/xwNA/69MMdZqyGl9ybMa5ohNuEsyAlKz0DNHAYMcYHdPzTF5E+
izxuGBuTsss2rKO3rZaC8MmwKGCUvLeV3XEJ8KTRZA3lAih4DlzieVDGojL73kjGRbwqhr2lWSY6
83wKJGZ7vVLgt8iLs/QrK/jLEuzevK+Wgh2iUfd14RT+HCtEqPN8IBxl3M9tBkKiEZf2k8+QOLg0
+8AmfM1aaWyAS9OFdQXqzJlvwDmFp8K22NErtHp/7lMLrn8xB/wCTFr3+TkclZI0ifH+Gh1Dkaiw
RWZQcp/xS9/0mB9xquHnyOEP96ZThhsE4pJExo6yqfzUMElKTXpKGViBPypbkymQoaULMaI0+fGT
gGhCuNpz6OodQrSwO5iJCn2eJZJ9qgIGcBj/mTc8CacWrnGqv7czPbpkft8Of23016b0qkqud03E
WLl2LfTbCRA1Uui1PAbmAzmVqoJkrJxSibbsx80A8c1IQnrcKQiaUVFySTYID7Rr9wnQEq97Bwxj
0O8urauvF/FfSr83Huw44uUrGQH5If39I5jzdiG22onnep/qxz8c6zxsIadd459wknfrBU1DV561
KIZ4wy38qada1iTxNSHIDrkQgn1IEMD5wdaMJ12BtYMJ8IYmP/AoqEQz/fZ3OhqrIqXp6pRFkcrH
m15l9jDY14VsTvRLXPVuNOlLJRcLSxxyTX0IdrYqtt5L+oypDQJj4yA28bBgd6LXmHw6vL2twPDX
Jz9S779NLfa0OolgBqlRlL4ggmu+zWqd43bEUzE5J8lSez4C9zpnQuf+OKjs831x8JMuPNyAiFha
i1UtElX9ADraWDxT8Qii7QtT50BAvC6PBLYw1LRiYn0L8AfFdF+yhnJckTJTSCb4Q79eSJXVgXkN
Cpl3LVDRGlL6TcayZ9o7gDFwBFqYMuswlg5EKm6LxA8J2X813SzLxwWJEwcxmSLpzAdVUzxHUWOo
jMeE3hYzAIOoiyxzXz8pqvH0KNS9kyVnpaBbGQU+lZWp3rl0UMAiLnP1Yqsda+zzzvkvKzDQWZgQ
S4M+4CiCLl/ONBC22ux8YFRfTi+lUx218uRZtS0XV22OBR3be6piyDeakPIar0lzfCfF6vrGFa83
4ShQeQf2+G6IdPoTVa1soZtytRPcxHh/m60ehppyN+8sdQXbbfO1FYNMZwQ6GmooiwMl0GN3KyTf
kWJ2meJVyezwNRxtNDJJdPLH8NuK/sdxaOeLF7z1YnTbcL/OYJrG+369Ga2QYrsPLnXghbEar01Z
S+H6qaemTLetV852xYk6igyUjwqu3ranNdQcLzm5U+RMHXVXWwZsVKvDnrvHNxdOWjrsKPuW+yJD
4a1PbCCiMubxtcphZ59NZYHp924cD6DDI3N9n7WjOD/yCx4M+UGyLHm0bJzmmXZ2P3cN9QLEFwcr
qC459H6l4fWAuVzymKqc+NtgT4KsCUVbNIdLZZkteYWRVp43KwbdpMI6++HBA3DobSDHjxzJEfW4
DNtDZRQKRbBSCibk8JH1hsypaszfF/IajzW3CfNwxXBcDj0I2HXgc/y+PUktnt38TIKdAmTtEHRU
vBVRM5vWeXhBd8gkushlazBGlJjyaIprI0b0qrIWmDROjspoQyNAYvXic2vRJ5nxk3zivfPaCaEn
AuDDWUaLi5kfqEwNdstV5I+69x6BMt6LyVAUsUJB8yOW87ehxMAlesB/JealNIB7Yl9csooQYXqT
S/+Jdz5BL3JhSzR78/nnJ/TTpaGF2F840gBLkAeu7wW+agvjW+R1mg0uWHNV5KqLHAiyH53mChaE
nOD80cKvLDaFsjRk9yCOeVM2HbMZI8YGjzVjbWdeD1/oqtTw/5jjNr8vgSGtEzciqthXU0WcDP30
2dbit29FOX1oBc1Y3SdZBuzMaU2K6LBXvtTYqiQJBEI1j7vorjDOeZNQ2aXI1GYQBXqIKSnNieUJ
eu09b1e5hMECOg6WuVmDPPCHp5RkvEe55CcPpNBnJH1LxdyP/EPEd2Vp11U6b3QjLsLGIdgKSKTq
W3l4IWIfusHdi4RsMxWfytDp/y1rWZQ9zHkLo0zIrmTklGjqa0vnVwrGHgw7zFJ6c4+AiPKmN9fl
Elmc9WOz+Jz4PWbrjZ/RNM/mizeYuzjfSHJAdiLN9gNQr/4ouC94jnXcG5I4EBk5BG1TR/DRqE2i
FNO6hbQIneO11zCLohcdjFF+ZdszDuAa31Irrfc3rtOoeXHaA/Wp0NCk02ZNx/RvQu0D1vxPpydj
tFPzES5uvtRbGywa7wKXM+nyfVHqmXH/xpS5X7NZzRmdLP8xElxMuvSTB5k3QP40L+VC0tWvXvuv
ad9iWPnGkGyrixuuA6ccB36qpRPJyrh5Ufn4nwSrzubzOx5YCUoP6uR3kLQDPgLDwwFisBM8Z0Fa
7C/nHRn+73u6i69Q5dHLn7LuBvk16yOs3O7X16vgGpAspAtU2jTDyc7yTtd9SEmSYeA+q8C7L2Yz
qZILdtIsLzWu1bNS09EEAHdCiG87UMCQlG99phpvhph4Ky6gZZ5LXyv74++NnIGr2GQFs6qS9fzG
llB1vsbK87V4kvEskA3xekyQRa9xIqBDztAw7x72R2t0uagkiucRKkIAXyofPtJQcXad8qMJLEtV
kgBrMj4JWCWgSR2dE/O2QvaGOKOkCjBu/NkWtubklpRPd9gJGD+rGRE57gUgTgVNW/xj4WP88MDG
VOE45vHxRmM+XjDiIE4Egx1xeIxyDzVD7HwhM4PydmkvYxjKvU8Q2L265M32qVbK17gGfgGThg/Q
qHMFZv174cLG4WkEVQEhzOvengf67SDgT3ERwMEzCE8spa/fkQalt/o5/3q+GIXfMs5N2hIkt+N9
AyQKpuGEmcPrwbnTrfCnyRW4H0TRefKnVugjuIQoS2xGRoIrS1xAXSZaHE2yl3U+Fnxvtwp9wr4m
lXJ4dkWqrka90xMWmQhSJ4wVBFVQtReJyMHD+EyFN6/Fxpd2PY3oTNvp8semnXAg
`protect end_protected
