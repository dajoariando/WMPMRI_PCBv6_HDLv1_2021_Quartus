-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
gyxS0Nn1rJNj36oMEWrS0ahuau8N+OuV3H808z/meqeqQcHAwE3xSL/iHoO7HmDWs2xHn06v/suD
HYwEG9Lfqg31wgOEsVZ7zoJF3PoiNdU9D6YLpWypWtwGji4hr9USAI/X4RSeOTawFg49CoVVq67y
J9kEcIr0VdB6Nfp32XIYOZLzxh4D0V2s/tj/2IjLnEC0BPVfH3nV6i5tnurE5j5X4ZVgBFfMoYoc
e4gWP/HyEiMMFNqQxIUsgCVWXYi3snywshSK3q6WrsVzhQvO3UMY/tIqIBL1QDmRMnvACMcGp0Uz
tiXneapo35BJdm3Mjc3TwYYlVlBgMTqtuAqcLw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 24768)
`protect data_block
maD/4TcSZRuqSf+78VmVAs6gj7imd1sR0sZ7cXKQeMcAnETBB64XrJOR3drrqFaUJi+fThTOL5F3
KnCFjBse932SSU6AyRrKKKi5mdjnsLY2x0C1IJKXrccdTMmjwCIZ5qaKnCZnPY0zGWLjjhjjAoGv
LTNgXe1rAaJ0G19WqCVBxVDW9rTwwp1xhTlftncxXPQZlo7QRzrZRBWopVDYceG+ixtrn9KZArBG
rMm15Boty0+xQhvv8LccyZGWsRTezBrKcYEw2PgEnXQwpsZgAG0TH/5b3CRV9p6zJsjJiMjCDEVM
DAXUeqrVq9GrN+N7TBIN4zdSs6OSGqqa1KVVemd6d79i0sSuT5J8eUBImOCXKgpCaLCd5keSGQhV
kO6tTNGqHWCiPkYk3zqBD1YGEQCPOJK7PW4KKno38h4gaTUhqcxI9wEFpQwIyfXCQZt4tem6+fMR
l0fS87MJNX4Ef6MqOLiySH5Qrf9C8r4CWjCtmWf7QuxwULjYesuP/quzD119bByINo0YE3URQbki
jkUgWpJktiqDfp8DSC0JwlgRioJeb5Nf6crNL7eiLExAdqzHHsTZYO2ctfMCBLQ6i1TwyJg0CDbJ
vRmhBlkOQSFCEGUnxEsh6CNksDdcuSDJpS/FxviAalR6otwiUo1kcFUj/srdQDQFSyKm+YUskAM1
ytK5NL2RcluVwHY2PmMKG6UJTlFLC5NqyDSFOMF1+a+kiLWt58tGut+V2SpS3AvvnfMlRLMn49Qg
mQEDAtZM+pI80Z23LxQXKQJfAl3t2cTEzaPTUI7DGMOXX5hE2n40xXsVijpsmEKcHhdycN/Qqv05
8v+oUv4jCHXDdxpw/DQ0AKvXNjJCrCi2SPRr2ytlipr8oe1E36wHZriPmeE05x/8rjVNiNmUdI61
Waalao75qGHAk33mB+kMWsl4+4BURDDTpveKM1Ooyq5xQJkUPg+U1c6Mc8tv3D20LycbfDWfb16S
+zzkCF44zv+ZVqqIStKs/WJPzalOtQDadbSpB49tYWHH7/FYz4R4rlaKjeHflAR5enKAUnjTRmLy
Q3m20S91UMUdWz1O4fAQLJxvFhsxyPw/5Lo0SktMzndMz4S2RcZ/wb7UergAVOySHAOk+Hor49TH
1kf7lUcWWh8s8AEfcDEpjcULFq0+0SpVcbD57eCaszft4ghYDqTp8WmJTBaN9pWnFiEQFz0lXEcb
x+5Y8rr26iMVzyQIMpDHU2X53QyUtYtLDgEQQFitFXHV0ZOx42NkMogyLziZFLPf8/uWnJRE7gRD
d/S1M5hJKJn2d6zY3vKq/9q61zcWYQOO1p8EudlNrEBzgJbtVyVGJhX/oil4wxkb3DnqFSVlbXoM
DnjfAiJQKbHqK8MyzWI/YFGvaZhyGP9E7jh6fotckkj13GBjVnMeCtLbvd+umXdtEzQP3mQwS0q9
tadUmpCD2Ebdk8mftSIZaH1t4bA5PyaddG+ALtih8rPJqu0rnRAtsqpaMlamOK8CuJSxQogI7udm
kB5HVjDeU6SQShtglOhqzOSR7Yz7e/C3rW9Z6L3rgYbuWzweRQJQwqok2iq8eJKPsPm01h7LD0NU
p4kjFeDh4NSemxH4SO9qiNMgWQtAMiyAJTTh65MbH04eO42UGTGxlNTokMd/PUbyOMGgFL+bcnJl
J1L69yp4iim0mVrnbPWiYOb62SH1ymTAMYUVa6f3N4nmQtSHNnCny6LCeXTggb+m+0eH6aG4Ln3K
eYTt+mVuS4TQm5A7As3ZCzHFAkVR43eB9XRweCV+zCD5IuyMMC9CrwVPpp7TB52pmwnt8kxm/6e6
acrICa/pD3ovQuWvlEEx6YuLk7MODgbJuXqJeOeyk4n4RFIZF+t1uYtpBz1+Y78WmlHxJvyQ0mqP
IhHmOEvUiqDCZVFVhuY30RC3mquiQLf8+h1WwygDd8oiSeF4SPPfrYMU6b3dTnZuKxx87wA01Duq
eWCA/T7ZENKUjQYDdFWgBZIq6T6Ug48v9txEkyevNH1skNHad6s/Hogr1MLykp5joDFBQaMbVOVG
ktU29dGvaAO1ob2d2dqZx/oS5GrJnriiqmzhhibob0gasic3rUzAzBIFByciu8MYPUu1QTQ7Gp5f
1d7D+OKzdVghP5jAsJTR2f+EkndVqbFS8O1grvaynkCxQ19G3I1LfWy+DhV/Yce3gSMdCom0AvyT
qUaP7ENJ9mk1judGYsYggekL8YLVAIDNErAS7AAcKUzlx1tog8vuPNV4D5OEMqlFHnW/EEb+b2Zo
+1fdXpUXR/bab8exgxybLrq8X2FndR0lj5ohBIK8gRmu96RmJ+mch5/DGkuMeyxZOjllu2pYsHub
kG5UdGU4tCNujpS+D9GFgXdxjbpsxHfpdwugqgoxoM1ZrY+AwW7Pzyht3syvSY2uxawjZWgUeUUB
RsmXK7+kInYjB5dRZIjtO8Cw4zmu7nV1SjK1osSBJfPlCNso0JRP+C46fiq08oPyI1COfsC1TcaX
Fc0Vz6JLTGdxyfeQabW4clmUVh5atKSIctnMUgayml1IA/9+4+bXhFLlJICEPQ1hkHbgFexes9UN
y/qYu24L8DuKox+EaKLBgy+OBJqgtvggg4N7i+8Kx97bwbYlIPLYZ+Gb58u9eeim/wOZjyGhXn36
B6EelW5Qe6DJcjkrlNDv7fQ/5xineSFBC2ZEZgr9zX3JnaixWnc3ZvBIFqTLL6ReQlf0MXWESmCo
1sK10ey8+/WrTtJjTThGI7kh7QGKZlzJj7gxAfPnQp9rx1SWjEJfIX59rAo70L2Qr4B51wdR853s
29W6TDLG+BemmZ1WaLPh/ITfHyxsOyXSROSOlHl1QPZuiqDwWcmU1YWQgFG5s1tmjm1g1sZlw8QQ
f0QtjrK5VGw5Y9oXcNsarN7zjv0hRN0aJU17cpFOrioIkVfOQFg+DqF2RfVP9uLbnHi0Z40uK9WQ
7/gRU2c4M9OLTscoqZ0C1hMnYNKo5HKGcHHeT9K9myj32GNrIJr40cUupwf5ZmYmrXbVXF82uFNp
1dJMMzjBm0hslX9jGMLeJmOJt7x7BphJ8/H8r6dOrQJaNF3epvPkcR6m5Mz9q02BtQvNqN8Ht1xN
pWXG/cIJenXbIqbftu5LxSUh7p+ECjq7zS2X33c0idUImgenQcW6j6fLYUwZKQurTuMeCDQR59yi
ueYh7/vmjoP9nAbkMAzCVCxl7ENxjD6cFjI+QC10cu14HLMQ/qo/eyRWj0b8nMYzww/544VGWtSD
JfC0bOMMp2Djxh+ktRcHR8L9JJtMkWthKduRnOizuEyVyGrPkzycFFIsEoM2kjquRwYasPUmXPA2
uKaI2HKLGVn9nLv8QtETMb/qgQDkrUwoYpbh2+ZYemkyhPJoUJhHPBlQiHzz0RNnouR2B19c0S92
mrUuYaiKwTV7QNBza4kZAhQLWtRW3sKPDKolDyhb9gP7uOK3okdR49vCzkB6R6f9MG8m+beqHmmO
lrjJUris/BzrrSb8Z81owqD8FfdjpInQh58W9BUbXZ+ZuxlvwOMzeRxMEcrbGFXslF894Fktp1QB
6yhvBxz5YCdOTzUbuhKi6tCzlCPS6k3QmSE7Mqyk5AjyXbCFGNsADj5K7yb3liao28aTnmzDmXdU
nMKowZUnkbMMtOfVbT+LKRDEvdVgXS9KidJD5dw7y43c2kN/jfwc9x0VS6D530W4We8A8I/8mAKT
mnDxkGC2neHqrtbHJMd5ZnausLoH5eYkEivGKyfzsc2hXDx3M3gZwsydVDZfjHnGNA2fm3QMww84
P7YrArWs1eQnheZqOrxNlKqckKw+QlbamKjLXT2IDAgQBdbjV1KFsXly50qtSFIdootPDl98TqqP
EIEFD6+d+GNAKkLVr805sN7cKx5EzAQ9t4OIS/uPYrGmmPQzxGsvx/q1+4xCO1hhXqoVD0TkxkVX
Mc4i8+85wrmk8gfTp/hLCB4h2OAF5ZEedfE5h21PiTvfUPjQwBB4bN1JzpntvO/44+T+ipct7pMH
KV/NixWsOjf5wCLhgIj9KSkQ7On83s7IB8tKvYqwlOOfvMgWY2cZuEepog/9jiBwozoPandESqfc
xKIWK9lXF9QcG+XOEKjCarZ4br9xNcuraZjOV3Ts0bnWgFqqHajW51zebDDyfvlbC95YnNSOxt9m
vE7F0LoA7dRFAckPNzfpu7MnZkBiLc9Bqy8RWWCVR9QV8ER1bGuwe9G9EpxOP0rH3EMWc6hTJB74
qSyoeGnwz8H2rST9ZCaGMjE2UEzx4ENztAS1/dBxO2ZXn6/8p46m83DOFFMuelF3ikNX2UWov4n3
YPHSAGvFRhTTZrfDX0FfA0AlYS3FJ+QpERXKBOBrmJR6HaDCx1f0F5dJet7GHYs+mSYHrNgeA7TA
+FpEF8tXNoUYZ5Oo2u54nWaaouKJFSGlAU2EmwY2jJKdAmS6QhloA+dVL0W7K+CudY84y2cgW7EC
LpO6jzjC0ZLLw6RK1DoAquHN+2e80nQ4Ju/cE4tZmjhhRfdvKWhzhkefHd0ScMQn/NC0mt7o0FcF
8U9ZcNy6U9hoDOAYXWEYuIy9P3r3tKnnQo/H5MwPz8i+/TBC1zh0HDngj7OLr2aR7CBxOxOzSitH
5y2QVnu1NEkKUbtgR/KOsg4+8j4moTiRJ0RyTxihmC08+cXWHXOmXZqYHY7Sq4BBV0eMk97jkbSw
j9s+rGt9J5kyLjXzCUmACqLOOrAU0KYgiHmbG4hXw994+FFgJFD/8wm/gkxt+ok5hTKTBoWzm5PE
+khca8DyY1T68eJabR2nJZc7YN6EB6Zb/cKv3w3NEvHi55lx+vHC1TR/6nevsku8ZTCMasxkhqzB
r4bcrOGwm3rupTPhkqII9wNAtCmmFkoZzfS1D/rwPsiLEVK9BQxKxw1VA5WWzmkfu7jbGGzSn5/Y
7Ww1UE+ZJsPLNBH2gTloym6vVkcV6DecA/cXhEyEWDBgSkrgs9mvoGJSalvxOLF6C0ePeNAUb0VW
Uh8J8gLKQmPeEN78IJpTFS1GsuC2WGerp8iHl2yH0eSMU8XZo6hz2+MSG2iVoVJsTOsC4n5uUsBW
E5Yf33C4yOxmFokz7sur4kgtSHV7gBf21diG5gFEfRcBV1lJe+stqEVW8B9eWFoHeuVLNOf3zzT7
kXPp7mcfkXCuxNWJFRDZnbxyYMLG2yr5AJo2p+s2MDpQYhrxz0zUA8nPBOG9yHUGYv0VZpLyxELA
5fbD7RnSBTduMNED33b0mgcpVvsEsRPIIykyIgUD8opGonxfTI2BXzuHLGOk/I7Ra8c9ZU2J8Tvy
ViO3oaGuDfNq7DjpZS5itAJypqH0LSoaGP5MnxQuamdK9vmMxEve1sGk39ojrqKfmQ1J27TAw+QY
uvQUi2NjJjVnTiOegn5p6ZcrXH5O5bODQz7IvidnTpGSZ5Fos07aM7uKu+BpEBo30nxS8QLx8+f6
USLXvk4xiy9eFg05ncl0V52Sb4wN38wWOX2zbY9FFVQ1SY7ZUSBwyLdl6oOEav2hiY/gVJaQxagR
65l4O8SP/Fng3ZK9x+7Q5PfbOzaEffxWVU7oRcABOuhuJsugv9jNw8HtD8zHO330vkK1l6oI/nnk
k0YLcsLO97vsxktNLgnCIjkoyxkzSY7hYXzoCXS4FTXbGZ83M4gy2BryfRpjjVhsitNoVSy5JuGa
iP6IaeUj1XMTCREZhBpLinR0N/E7CnPfJZCFGGLV1dQQ0SGN4hg6T6SHjwPakE9bC4EO5zs3oMRR
L36ZxANkxpS9W1S/aoolk8sDW+Fu4IboKVWY9wEDMIAFfxB8ghxvgTRROYS3gsQLhkObi6ONegSf
+U5/AAcrsheLcUiUbnn+raXmO2e/dfUl4pmueF6k7JnrigLuqw+a1Y3c/HgERWZxd2U4YSPiJCFp
05kSKIybIJjB8RYWeC2u2tUpYQrvkMWT2GuDfDeeW4DKOaQCokJxVtb0vC9kqb0OCLEcadxPdMGN
rkrmoktRcBewbqP9HDnx5f3PU50wDy8QzdI0r/Y9Yun4jKXCt1VFcvhH9wSoHlpQsrURUivF7zcD
t71nCPerdufw+UPTLwtTngtxLiTges1BC4T12xND166HvXXhdCihtLHVRtceszLYZUnrzz9VddtV
Yb/uTb7n0skrNdMEaUaGSgW1cewyF1VvT2flW6692/BapdVjEtbQ2TkedBBCwOaUKMPrCoM92X9o
E6xMdhywJH2vttJPQpOCy1QXaOoJFAxxR07J55vcKjx7xd3QZEEmm+NrZP0yJKIOxNI0SPKNm1WX
jZXkkwnYLHfRI+meQRNXt9onvqk1VwAgdCob+0jhwklDo8BLs0YNRZY9jHHKz703BdULoFUqhE8y
k5M2WSSjeD/5vdnOzHjhNZgUgkALibG/H5O8ngcq/8WjCN1RS65UodouU4gRt+qSA1t9UGfLvA46
VWQyfYVCBJ3jrADdjGoIVfTji2BPULoiWqffPWjq06O4y7H6Gaqv4mfovKrcL7VJ52DVhNqftBE9
UVwJS6grj1XKcxn31vN6dRsdVXfNl/4GSE+FPxJi9WW3D4dJ1pKgTNSkHK0QJjJtyfDqtDUGfcGW
or18zzyVS063D3HVYot3RcHe9LWNmK+8yS91DQb9dc9+43sb+DpeIJch9GARoo6kkjly+9QiTWoe
Dcdvw272qSJc+48TwRQvCGDhpkfHCF4K3P3r+1QIkyRrY6Q5BO0trPu3YvYK1qZEGdsEEVcZRrBT
2Fcq2MTUrLoR4K+EHqCIX/146jlotFQf8w9ihvPNmlZ9FM8vw8ZKPmQisroodiFvNmXe3Y79VRFs
ONXvj8RjdKRGQGDhKGQN4mpnVtJasSsexk7ZGDaSmartKavQyas73jf6/+VXIbZvznXuHQQjAKlN
rl96ykuJXTacuI49zTArVZCV7R+QKukoWkE23lg9gp2haYGkhhhCmW0hO0knR28yVzuWbsDTd70l
AYzWIyzweONkAYyYpg/VI52gISE1mRdYkwI2RK+wBEd/pFIGRSinax+AKKeSkNYpl/eC/a1Lv3mN
xjgKVLM/1LzZo435x81MSfI++vRHh1Am7pGh0MlxYft7UlydnFxIPr4BUU9rWHVnaNhqI63pJKr8
hAF5Ou9z4ItIrQ3Tz2nXqlOmMVIdtUI7H89qS5gSLMtw5rvbnXWdfqCeVPC2t2VwYdkqldT/EzoS
L6/E8XF5kau/Uqd1yEkeZOjatxdo95d/jxTmQHC8YEJHouATsRNlG+pYmQCMGOWxIjT7rFuNiXr7
OTkhySzR8va6mlkQy98CTQNDu8pWW+spnuPxiRJXC/hOdRt0FTBLc1fM5G8NzvOYfRXtUnobOeyk
2o6vf3Y9+D1GIQQ/PSkuwo3i9t983PdjGnETO2F7tkupr9rsqxAj0Y5jE1c5SjpAEzotCBacQ1AK
RsGcvBFCiQPSgWXO4W9U5y6T0w7hNLXsYT8E6Q7NgeLYSsFOlxxNCO2ERlSu0vHDJGAMSIutPWGx
JBIcAxnGpfWYfDWDYbX/mZK2Ww817ik/C7UTwRUFL5znRvP6A9BO+9l36Bjd1tfJVVUUBHGj6GZS
CWsmC8ezP66C41OpTj46pQJO75Wz3OSeb2lGR/SXX//5cbG073oftaJDq7Uv5e8ango8T5QCVOWo
jgxOIzLCH94yUQSxwmJ2oP52Xus/Se3u6TyJWdYWN3bIqe0nI7XDgpa+CmXBxJe6imaKrxYTshJo
FMlAjUL6JT8gn7QkLYEhrcNImiegO0yHwyGhrInMzzswSjcADNRUSN4RKSORNyx8l7iPJaHgoIr8
Lda8HziINZTL3OY+dheqTnNlpNeembGZItyuy09Xpt+zyah/XrJty5Fr3Ix4VCLQrI+foSnsQF4o
w4H2MvA6Ch9ecxVLt9K3bxmMwqWtRivYaMuD43AsKUMsGBFc6qZl7Z3hisppVRSd/RA00/Hx+IvE
nA5w21yhWH0UrlUwfFDGfXaBt2arIAyrlbB+V0cAhwfs+ufFOfJNveP/vK+NhnJ73GCzvMVBYz80
1K6DwapkA2ODzgOkEGI12ZFF2EdXsf2+M8hLGbH6wEZaYZj+Nt3zas6g2TA26llHQ3rxh+1RbGpw
DwmxfcezxwEF3teQY6rX8IhzA9lxyAOl0q8Pex40NCHDCNPK/Un1zHS/W3yoHeworKnWu7KqinUs
O81OCVFo/VufcVtrGav41MNh6sLAMsJk1jbDJVOeG7vdLBOzO8/wtNB3Y1y21rLiOFgxt1Y0XPgA
66BHLEFbMK19E4KndcZZbErBqJqOQXySVz7BXIjqXQwlmkqVyEkAux0znW1ZSHTormxyDiJWNtTM
YMlEawbynpbiK70fCLNWVXfvRlW7obgV+WHudz/ElWkjyC6NEvCNzLV3uiawwFsic0K/BDKaOmKB
tFJnKUI2dseTY34F3DM6j41Hq/NPLPlOify86XPFfM8ccE22fAAnqoN70gDFGXJmp6aEcyM/NgxK
xKqJG/QGm5m9wV2pik53FCQ6sdng9vhdfvqRRRRjG4MQN8dUrTK31Y1/GPz7rJSfGQNQgh3o/xk5
ed7GrXtMWefm9J3VLtLep2nA1hLuxIaqHu3JoxVFf29DdvedN53ZJHiCk893+8ZGG96oXEg6JTEZ
3Wx9xVNEE32uL/7GiLiW8yqLK13AdMwUmiayMbaoCanTP2qhvdXIpt1+EZLwIJZdAjE1k4XWuShN
6VJvIU+J/feXwdhRRd4c4mtvNejWPitzKAM//8UdGdfFsU6I/6OPZwFhjy6WsEUgKAspQ2uCgJaX
y5mJPyDBdYbdMFZ6XGIgn8KYVj+13jwZz9JzhPu/iwVASzgB5WcYDxPA6FuiU27QECRURLEJeR84
CL1AqBzFqRlT/Go/Gz/CqsgQSY+1H6CQD3BlJN2p1JOfF1WnMqBcV48AFb6SMXJlm10zIf9B092w
0Fzyvd+X6oekwA6WZD1s2N4ngPmHOCdJOUyJNEE0KmWWyWPcs55Plp3rvJqoCZ264RLrNCI2AA2g
WSNQrPNwuGzdX2WGAwe5+0L9Dz1GEyJvTaXVz/ZV+dkZw6POWXS4BXZ5LmUhx5WX2K6IEGgM8Wkn
94/FMGreqzrqNpQTJerzFQ364WOWt1cOvCS1osD7BYaOGwku9y2k3DhqZFmYOmTeYZAueQ39Kg7e
slDwB3qhfRZ8RR6EPPrH9RB+tkYy5QQOCVc4Gebr5tlZrDxVKwEgAybCo8eStWIYBlXQLPzDoRxG
lOjDnzQrhsxDafKE/EhwZTHc96NhX5rGEeUIvkPb3YMCvDuzdliPbCGNsw1/h3iwsu1vsxYsL3ma
53niJSN7zARx0Uk+YWsu3Oh8XjjI3MMab3FWTXP7GLyh/QEUnFjk/KxUZMXz25E+7EV2Q784K+lj
+6H0HhypTmenbWmKxNtrQ1K/AtvN/oCQNgMSKktPHH/0X6XJfGCtBWii/Q+5h9GFnhx7gO3h8E7Y
jk4f6uC1NmVSU+XLZTOUYNJyv6th/m/hOs+Z6wZDIWzstMVsh5QzE6gUF2NzB9UUa5ExI2MA+wjT
sLdBRck3HYMFT30dltQ+OqlQi072kGQWmixog14DsVJZd45c19EB/ftKRfKz8k++EVEwPZ0vVSGx
4l2A7zxDII3+qWYwDykKiFyaN6xa6cZha6Sg94dnuFHbjXrwxilMECABj3IQyNJu/svabJh3LiOG
jUHeRx4QOEo6eUpDvmLCOtSN+gAqueiF0+gL3mbengQwiAdYkOkTbWj9YxhUpW5Z+YTy1dEpauzJ
hjeMQ07t+PAYt0LgSkkTN6fO0P4438NwqcfB715b4V+bcxA7lcz+jcu0iEi7l8+Bb7aVFirRlrd1
OSTC7PmK85aXpyZ42i4iiLOsnMf9wd3609tk+vHQ74v1o0D9rpHRsGwPUci1G4oBmef6tC3u5Bfe
Kc1hTHA3bbf+DGJNU8ybDOWFhuhagfcIqCwx3lOdNmMESF9jsjJxURAEg7TUfwdQTcVRtidF3uz4
CO7xRLzPOow/TlwCB/y9SC+mVc5cKPlsU5sjGNqOxiS1erYlfembLFJo7Q1cWa8qwEwoq6FCeNTW
RpKHFNMGjygMiKbVRVKYJ5VvA8tRcQk2WS+uT8vRDavknq1JyzMCd0ZNsAzySeeChS70PwRhrpm2
30g7ABOIRm/NjZFYQT18dqA42IzJ6NxspccDReL4cZ9Ns6tePD8PeJ1OM+C7aDTXGnBIwFc82JQw
TGAo5zh4FC00a+sI8x2PExLEDOUJh2qkg6VPV9hqeJUWjOAGZ2pDCAQ3NW8ZY3vOzqhqQNGpR6+A
icsEmxVzsTDue0jXkUj2rMIQVq9qPZHrlFR/O4XXePsAgsafvpNxAepriE+SQOgOFuqqkaJBv85R
NOr2Wmop8+Q3kRoXHXv19GXB8D+rvAhCh+J0zK7wxeFJD1RNwoZ8xYgTRBLOkqpdpLZyrf5+Vi2O
vFKTBi4LaMaM2BdIzCENP8N7fzVzNRGMS0athrtOtJxHWYdk1x8mGl83ptqfNiwAx0hWn3JQtQYW
N6xAI7O7Zn2uqae6tc+pf0ILmQn8K5hXxAboX/dwMip95oQblDhy9AYK38KJ6m4OaXsKyVDFcDCm
heMJZJCoSf2DUtGS1YfcSNMLe9x7aKt/GKQzd6cqQ2k0ucPVQaEe5kMPpD73JluQM10UUIlI6go1
ed/ZK5J3ABY6WV9x77YLQ0IVcThwMyZtmcS7Ozzsj+v63UEAexOIf/0jQaKElA7okTr+iRuNv9jJ
U8V9cQDpVV5cZCILgTgdR48AeXt54jUh7Aq4wlL9zEMKju496NV28CrNGzq9aCtfZpsP5mvekLUx
50f+/nejyDR0q9EAGnpFVSJC9JDICevN9vfCgRBEXGRwZF8RM3ybj1qjKqEdS7Y+nanCLqbt6RR4
i3C/w7JAlDHX4ot1/ly4OsIFHTlGn54s199rW4j1kAnkEwD51Xx/vv3qrug00tS1HzaXkdP94qSu
Xhmbf7PFR6lfeu+owwJzZ2SPPUEB/Xrr9oSpxElQNIlh7l0F6agXGlvpnwxJjEX7ltQvRuyMqkBZ
xgSTCbrAYU1clcfdGgvEVBENDT9jNZtrb0mImBPqkZOGgHyRXGRYJGXG/eG4lDc3nyfdH3+NyYoZ
TqJV+nGwjwQ572+bMDdAX1Sb9DUEKN5DOgwpkEMSxr2nSIa+EB1vASFsZZ7Ol/V8Kzjhg8uXEi7f
CA7P0lkLDim7wGmMHSRZvqJy7pBawisUMl0RYXVIqPe5MuVCm8HibFdkSlSEp0M/EDSzeifn6fcT
mQl09DV2gIEESXY2N4NC+oCT/RhXtLT8v1VeVSVgdMFhrgl2E5cIHS7iw0OVjuQVL/9yIGHFWcNd
qBka+uYfA0Rc4uceCdWLoRhBOYS0glskQQEqdmVPlLpRtE1E/VqH2uyGIj73XbFzqhIgxMD2WaBR
DZI5exMlUpA4Rjapqs4NHl4Z+N2F+46BcWd8tcJ5afIxloioxtpB4Hv6enRI/XOZLqWAOqOp/5zI
1ERmSIx7O4kVJGG1LlfYeofzX3jWqv5oVC0qOCOT+I+YKiJCsd5+XOuaDZ3kebyXhoMjMabwsOmq
M73/Qn5I/ijpXvoDhcSEm1QsdJDrRpH2rJTizMkP6xEuTQfIMv/M3Zg1kSPdAIqwL0/S1LH0b5NE
Ix8SxZr/F1I2bGAP0EU8iTqySM/wCgUJHK+Woeb2ri9WuwIzwjXbZs43FSx9KuKkpUad8OcxC2dU
KPB6YItyjK1cpy5ypMU9c7q6DgrwIQXBO6MQhgBgIlL0lEGhaQJq1MKS4XQkPmK6maoRaJqOJBKJ
ZCh0W44gVX3FbXDX81aMH1sV8ZuLcKJFQ4Cc23eUMlbemnFV0gN1PWe7Sei+qwBKjv8gvgF+B+xy
COev+u7Ni3VsAFo7W0jt7xdNEWE2ilGvLfS+BiV6FtXrCUyO8AkKlVY+bku6+qmcHkaPoiPMSadr
Ut+JApQDNWah4VTNp6PIaKr1Hov+zAqzOGt8o3kwuTY3U+Kj1l1YtZVFrlOIGQe9IFO590d5QpEa
lF4+mzg3xS+lskh4NFUvgsTdTASyBt5z4RPtEjV0YXDaplm5Wwc1L60fHypo9/z+FlOy9CGvipQh
l3lzta9MbE8xRrXAwBhy8cngXOitMiuH91Y0DS8leXTzHWtprUraIcHiXIKkUEG+gUCQGHVCn0dq
XycL9/PtDsXQnplejPB99PiCuHl4920rCeEyBYBU2w/2KhoGCzWvNJTq3EifWDtWOmcnWC7u7EYv
9hkx4u5XIAtBsfQ4h5ya/N46snzMB8UwqEqDTA0W51Vtylw30Er5ReYrk8K2o2KdUYG9GcIIljsw
uJHrhp3Y1JqDXEZQhrjdQY5LIxtYfHDKoUYCha3NWVK0hm3nxZmNjWIgVVJXB0PtL02DOF4dhuYq
I1FYaaDlqdMWkb16roNVLbPjXz1KKhd8uV9q6yRfx5YezCrMwz5brGhrn1wCOL9wT5VUuQQiKGic
3qZWWL/Pan7RrWU4OFyouGLCusJ4/pavfsEL1yvaFwydL/aL/8qQ3IPOXmRq65iGzhfA713Cl7Ad
uG7ZKOUoXy70c4d/zn6maNUiH3SyJTWwXBUU8Jb9hHHTAaU/uXh0nidg1nkUuSaHt6y/E15gHN/o
FcmYI9tWamrEgw03UvP1ZSnahIYT2lslVIz1oK7zuTC8MQREE9YvGhmi+5+cSUON1hbMryM6POq5
umnayTUPKsGX4svUkXZlR6adKimLZfrWn1v8AVHfAlVimh9HguXAr7fe3jTOLoqNkit9CAvUKKk6
yssKrh4bjloeAjESWX8C+owksBE5L13JurdqG00DeLgRKig/SMiZHCOfKrKvRv1wzOyekhnfvMpE
lbIc2vfz8IoL54W4OB808mNZC0K+x3QGzHcKNf3Zghjw5+ttQCxUgBaHsbrwWB44k/4sz3rJmAg8
xKRFdPSw1fQdG5ZyLzCakqsPB0AoAYUC78oG2pbn8L4T3wq5OBypLzIec/j7T0TIwTmQ2Y/+ri+q
bSJH4W8embD3UdGfRhrWfajl7RmnjPs7RhvVnoApsC1Nquam65RYjQIB+dfzBqxGj56BXgPwvme+
H9xx4oc01LtjD5vzODFHZITgzKsomuRgt8+VqN+ryU1qBixmgUZPcNbE3NvdvAtDPsc+90NE7YB0
jHlfK1sQxkakI2iOe9bfD/rrtj56YiZze5sixKUB3LU25z94SXsZj1IMJYMq807EKe9OBCOy2xwu
U8Vs/AY/KdqL5cIVsrfu0XTiQbhDIpE9QZmUuMTdU7Oof/zS/PVuZESSdjLmNjsrUyq90ozO+h7I
mfmOceF1fKmPeW1yBvehhu1GeNaChEVPQmVCRah+ykQPqR56bQxU898ZTsVEclMuIviy+8Cfldzl
ytdd/zGxiZ0cRnPteEdGBW3StWS/vQR87rf5q064I3fZzqjD08RTFaCigsrCqq4xLsWenMum9NAb
762w+a4Nnkk7WlsFInOS7Xj1e4Cn0jeU38mgiNjdd13P3T4o2xWes8vLdTo35z0OBLtDl1+zoiMj
R/IloOYfGPOHTpP6GYvPP+m2AYzjpFWz8+ZzyZxv77AWcIn7G7Ip2GkppyGUabT169nazqXbB4Qk
13IE58wp+GOPdJ6/2pY+k1CO6VQcrDbD1SeZPCFpEbMGvGDAa4Ta/NBFsjzb2YIJ88qCwWosk+Qf
OBCdI10PmHlR+oPGO72mbYBbkOYHqhnp1qzUvGTTkF+efWmHlW1VhDfqvBymDPkufoU1w0+Kgp7M
gz5HGMI7xQ3H5c58IkB0mQPCE8jq0S+3cPSzwFjTb8BMRdw2DsTcOT53XN2BLvYZldOxlpIgEB7/
4CU3RspTGG79NnKRcw+9e9KOHJfaNcD67CtqcFdnjXBmlZID6c28IymmB4R6FqW8TIHrXZUhF53Q
LMXpifGJHGZmkmR3QeqwLmbPvrr/hMdkCt57DXLKd8T4ITnGPpAnWwGkQS3uyxq1eeYZH8f7RBer
uoHjx2Nlv2SIg66+NLGuwElECb08BDo8MPVwYNTteG5tTlh93QjktI7wA0rtyNN/xxSFM3tWSHs5
Fh/vtAGtpGECOARlvUA429Kg1h9JVx8k794h/UUFeiv6Sp8xOMYNqueyaDQFXSE6EWTWqSFa5y43
aqF7hg6ABhgZAeQXaVDeEeuKtYZt0f7gRbKp9NnrDXAoI11VARxrh9ZGTjxtq/13I6GIYp0EEdkc
gsYuxVKHtPT7F8abEZEFlOE3lolH5KMd1JM3pA6HwJapuIdoT/WSVF6hfI8EGY0IVpvC0uGH3dp9
/94Q6MyrxgSZnDHiYqUOI02oujiyD7orZ18rq3fhRr6A/OObyqkoGf9X9O/vFUuxdgYbH578xcjf
SMZYDWMcSFL6SNz/DRiBWLb8jshgosCx1morI7vDuN31/lEaAUBgNKthYSTXjpZjvHvYaiuuAVxG
Z1Kef0aftdPefND8hV07BqEq/B/7Sdtrdj6r6qFyzYIHVfQ4DMc6m7wnW09wF2g49q+w8Kd6E6NT
75O3Y9/7FNv+NUEPmOv6oc8g4P94yj5+3Uj9rXWKGBnpXNnlZs8+Ldl+pRhn+pmfLGiCVS64f7rS
3tq34NN1uyAPwmMFG2w+uXxbefuyrzE3S7cScLImYsXv31UTPbaUpMRALt7m/hbnkKTz9pZyvE7b
HqSVj7qoK35zGBo/6miRi6CrjiEsBGFUzBVKktw4xl1J1EMWVyvx9ziS+kxZ2/j+8NGPj+fvcWGr
M+hgJTZm+lxLyUddSMsvpAa58wGN9ZYfUCu8fDCL6/TdyVaCakYrvOmx2ZZbWKj99tJ9btstkbLc
wyEyqkRnD4F2BuAR5rWg1cWW+iLny6fqCaiJcfiIZV5okshZbBCQnsdSpzXsGR9c4YYZnTmZ5K5P
d1XQM8QPdAuxeQNzWbV/IAV/fjX/jk1ZEhtNT5JCb+uA89YGkAmKytAhvl7FDzsfVKz9SX9SiuRw
9y6SPQZV8c6GOUofva5D6I4x6/k8EPkGLQzgNFyjA0MLtXbDfjWuTxGDprToBpfkBJRKVo18ykwV
cdZgb+0SIHvlu2ixc5LsGXXbD1sWfWmbUQ875tJJoiS1PbRQsCmXQUmjVgrEuEWjn+LyqHkECwJR
hpMHdCCtNorKuyRY1oxvQLcpg2OAowhnVy9qU4PPTBiTFlwxz7sMrv5AkJ8pOVgLqVoibJgnGlMe
6OF/W7vlv3qj4D7+eok8nK6CzTZXNPIhUgH4IuULoFi6cnQxWs6RYvKz6RW7O3duwWAN9ZEaDICP
44vAM80UjkhAsTN5WCrPbLKAmi2qGIITBQnAOY+qMRjHer2yaGOXzgBGm2LdCTe0j76FavbFUn3A
qlp4XUHK/DT+3mCG8dFQtBCNdC+mKlk8cdQhH/qWgTBUfTcHXAjQOswz4vhB67P2A3tY5vmpQ7CJ
xBA1xHcEmYHVEf1ak38P57N0OtWxDk60weSkOdr8aBPFqhFJGTBFQjAIfwcYdijkrZbxfTOR6pgE
54otnMnG7Mii/BqLOv+G4OI5Kl1eoNFpVCf1RHWcu28A+G1EsOqKyl3jlpADeYu44vzKx093LyCG
F2KQvi8whyjtlpWgGApcHqQR95os7jOSofQ7ygjZK+d+Y/+Lt4LyEC7T8dGAffc4RVPUGqeQFpwu
4A3VWBHZvcwe56v6SsrCL/P/3uv9aBWjfx4raUNYXf1W+IM1NWjuqlyL4Hc6kChpGkm7U9heiSSF
y2Wr6NV4wrVco4AKwq1LyVihAD1Pe0u9M2iUI1/pwdz2mrkOb2yywGgeqenNyTxrfe5d4Ws0rs5X
O4CbkcxmpVchqtVu7phLdkolLkIjzDo88w9n/2GtDkNVbFc41R+3kf2lNWbLvG+n7mNx3+ECN79p
qKodhAj2oKntAqhOoyGVCVTBAKQKxlb2UibSSsvOFJmMZWjnfjVLoi3BUnuwaFiROr2QWyLJfH7v
bz2RwHmYOl9TA2m/MDe2SnKER6HOB+o4nyoN40V0aA8kLffTb5kxUzYm6YCLZuzYoZVlIDeR7DJV
fcBfr0KqGX4kdDRFYpzIBJ37FKBn0yRHWWhVBzu5OM89qtgIKRvzAQYTnAVtt5XhfLJLOu2u15Qo
o4HnGKmyHnK9ETcgJQyMhIt20x5XrFREEkGAHR09KAg3HuhVtYv+mNe2rD26DlzudKVgj+S+JKAt
5H1fUkdini8F/pumYOsLdf3j4vUlmqdFUKS6691p8ooy3Odi0lUt/brGKSJ3Gsfqpa7kM62qDIW8
PXSukE3z8/v25MCjsmcpWC4v1ngac1mYvmIFFCQCb7C7+TPiKT103Zun4WgUE9s1dJ6ChSh/kihl
oyUszxVAu3TEGGK4+B/IcR484Ag0KU2wckfCNkrmEYLEXYUyMPY0Y7rJV6w09YJw6oQYaknxTEcV
AwKOfgLVXNDKKPwZC8Q4W1CHAbmzmI5vC2Cc4IGPiK36oc8W+yjYei3w2WD6vhwL/d5SKVpUlCOx
pcru0fXBbIHNtYWtZuxMtUjEbpibYl3Zc8zZP+uEDkgPuI5WVQB7NTtcG4e3V/LO0CIgj2TaCDEQ
GvROFa1jgGE0zR7wrO/rNgij9edAkqY3QSghWBgmQe/VNekRHQeuTbWh/m3QLrl5j4+5F+IigpaP
HEJth4xHh5MEYh9dRkD0VxkRF2fHacbjbmVeBKXRb3uCDrr9VL19O3uuRE9pvNWmg0gKSwLDOMct
XON1edJuaP7UrAPi9lkpxQX7lygwdIdXTGT/3B3OlQaGkv/iuTGvHbbqK21A/BCehoxf3TnwJrMF
OvtvHL7xEeUaL98/quzRJa2bEx3PxwKorDf3IInJiwgBySUecusimvdrQMgol3Xc+b2fwgeO+LTn
Wtqy08tHd80440E0Qma/bV8H9p37u+yF/ym77e5zmb9GdWJfhZbA7Y7pR6650tuS5vMYe52mCnIa
bGsE1ko1eQLNsAv8EdefhMtvuWed2RutrsrP8akXahwrwTdGh1/PTM0+VedYWZZ7B2nbD1apTx9/
Y3hdMHndF/dhN7ISMIaM83PlvVqUEFtFnzmEF8EwXNuHkJGQu07nFvPb1f2g1/lg93MpgigF2lg/
VeQoEQ6oBYEvu5eotZafqroTFuGs2qFDNKmjItfJWeLqRUzHfLE+lPecCFFgpox1QB07RN5rAO45
90s6oSXpAC0QyING+3hpJnbt8Zzs72bLGb0/LIXXIBWi2FLgszocoUQmwFTlZRbTTX2IInH0UAMs
u/8LCCUyZT4z6P78Y3yWyqCkPA4FKkiuOBd6N09DsjSGT1TexW6yfpx8QqrVI1DEaJpBW/vkjCcP
cFSIxY4q40lkyBXyimkyxuz0JiKEy34PUKflniAwrVfAOMgcbW/dssi1kO6nTYNBg3Kfn/+La3HH
imMUOItKL+xJx1NXl0IRTPxBGxVjx9OyZ/CctwetA/SyJsAlQ7KsYBdVi6JVF7Ua4ilf+IKjUaiV
HQ10tTbrOYIl8vAyFCYllV+CZEAofifNv13xJeQyMe936rTa4rUUte32fqAaBMtZoIhJ0HB05oQN
2mnHy9H5hS5hczCYeRuCeXNbZ+Lk0emKjQKmjeMQdC/4ZXKnMIBSSeKtKAds+Im15+XPO+9p6nWE
BPJDQza4zn+/40O6m/EOeMWe1I31dX4TuBbzeNi7zj9aSbYye3t5Xsp2rBHUGcXmEnrTWfl5k2Nr
fsG04g+7cEGg6GB9we+FPLE0EVKX/QKOge1vchDdUGJ6HaWJlG6mG+GQR5xBjhHtHuR5vFMdJo3u
mnbgNBL6k79hzg28pNui0XReL5ToNbtbr4mTRLSSuW6QpfTxCOMQB3b77aVF9T7MVuI0zh9zTEjc
8mtuKUIrsYIjDKoS77zxzgIApOWXLzdMwb3pget7e9IIpPzbB0jLYrnph6Xuy+cHDjhLA6W1yvRZ
f/6kVahWkk6m5uWofvE+yPJrIb8ypuICthADK9n0DzqYioeClLTuztU/GWXG1DAJjAckUSOIj0aA
tAaFzfxgrRXHJAjyDeyILHBCPiIGoffe8r8JulaBQb/oUYbDDC8a2vtA6hQRQk6EzX8Ny7KrcUxS
oNGsP511HGp282FyOQvccHnlwjrAZB4k2GLa8nNZ+idW4sfAZeUe8OXOnNUA3uZjMeeBuSyjgJnk
qntmTSJgn6cpVCz8OsIo0M+gi1rYa3vlNq6o4AjPTHb7mYkjg0HDB0jK+YdfCmGMq6chmezNRY/Q
9NhB0yhT0Vq5eY7N8h5AkMvQSN0PcsAnIHHjt6lNfIQAMkkfd0VrgGACXKTwG44iEbSYSn+danm/
NhU7HCb0rPpUxpnn4ADzxUKG5HNd+Sf9zlN+r/YlTUpMOYWpysM49t6+6zNi9lkBBu5n/PMbv7Tc
HmC/9g/vTlzyeMMEVWUediA1/HaLcKONa94Q7ae+21PSTGdD7MPJ0xscVCfDzSg4Sns7G91SwGio
L1fADiUDME2ACU4T/Gl8WbyxNgmiwTdI4iUWtayi31DGImDZv2sr+19kHxk4ERB7vdg6o64MYxJ6
rUgBPlGBE3gL2/SwrdFPqn3e15hyoP5AAmDVaGu05U3PlHb2V+tbijQ/VbL7zYcESkwb3lFxBV6L
0BukNEzmIgcpxBHQt4dQjZHqEI1qENcPS/6H3kXYv3R1rV/EsZkuKezDy5nAGURvQC5LVpXhlXVY
iZlJRpqfIUJ7kkfSVPuP6K/WEOk5WJFDtoJZ8BI/0WqKUytEZ84K8U+hXV42sNURtp2vgO7o7nTI
sVlpnHDXsC6Usv7IV0gyfyilXnFYGC1/C1bF6rrbSd1CHhPgKy5ll8SQmtc5evPKehlvIPaCDlNW
YNp85bUoqtxe4fmb8HBFBRC1alVZc8Z0sFX+e9ZV7xqzHrsbVbrNKc2l6kxK/eiPuIMjXGIVw5re
i8VU/QEMa3hGT35jhRv7Ox3KEwjhjrvAOJ4/clFPQ2dytayeoR6+3T3N9DE8OyORLs4DhlicZoPb
mrNuzVXpVRWmyg/rHDG8/a2ZnUSFC3py6D0eNtbau1d9gS6T5gMfEyk08nzJsf4Yy0+NuRTWLJUp
+GotA8lK25sC4aalqxYzvUMIpdgNMuIxD+BsHambEfO1rm79xFZKSobpJPh0gbgI4M75gEqRHRJ5
OMQdbQkpCfbzOtPs2kdBa0xiwnEMovLgLcJezXoDyDVKRQ8aXTQlg43tH1td9RG4SkxWWjB+Gi8R
xHf+MXVWdtJVJICvqcxMuusQqAtcYGl8/LOWTs8l6GwZaLv0Q24oiNEZFnKk9sPtPufUE1q/6vHJ
+SMd2iUx3gwNU+ta0I+38snkD0EHPfx9XP82jarNEIYvLm5C60f3oNRVCIMF6EFeTHINSaEYgm49
Kso+a0VuTx/tDHPKY85HhTCPfvXOVWBI7l2yqzm2pApKCk4FO28CKS/2t26AjRMSYQHufl/1tVYY
mdXlvUv/IaBMDyDUEZKIz5KMZYluiExkV2JRTdtwKx4fGyZFP0ezQxvU7lmDnjtAy9qFjVD0Hj/8
VdvcU8YQm+eEzNV8e00a4dHlo+NZWBecoAPj4bROSWyhfYF/3VKQ8DQKycHuGQnxlRc4Mr8Wpwco
DgaH/iMc0JOUyliVe3/WiL1WIBkZPZjiwUXdhue55pZ2Yh2SgDgSxdvpUkZi4PKK1YCYH6sJHdt7
Xmdqcb3oKzmz9044wbuCX+KSQc87ShX5bpRIFu4g7z9M7CI5XTyIS1erfJcwFfKlB3hx8gS5OilW
xKLkMFKj9pyQPaJ8iR9yLyYTzuNFKnhglBtZnGOoT68iPRrqf+IytKBogu5lDgNIHwxsApZYzSNA
Q9AEhTCcOBKJOS19CvRSu/4NkWzTLkGgx9mBue67elaMNtT9c4X9WAfeFmowALroa7YTiaFVyBCh
70CspbfJXfOi9NfVt2MJGiTzpnqbw6DyUf+HYhBUaPP5IzePlU/Sq6bwDLEGsU6S6Gljp83no72p
VZjHYGyvBBnxQMtr/Xv+yU6qsbGJYkNCzetXhuUg+10uGEjn97cmCYKXrm/I5dD93jnmPS9y4BQ+
M2MJp3+fJt0Hpq3jPyxz2SE0r5j6UkpTuSxEgHq5xERhy0S20jhYm6+a0s3T4w+GmCjsA5hFsXnQ
pzZ7AWyjmit5i8KoprlIYUFyyB9KzUEpIYRCzmqtmIkoNGe3httbxhhPR3fHarb91xUBnXMqi7fg
TRVzov/1zEbqTakQDn5+0gVyIw5aRO9zB5rSO62JXk/SmZBLv1vt6q87jnYBWTdByoNb1BfcQON3
N9txUnr1U8U4eMfw4m1Zmn5FuKsJmwpm+1S+SkpQTktRGKpIXMe6CIfCmx92GZVeXKxtaCMZN99Y
4TdQ7NFDAlxH4qjQGVh5AcWmio1p0lJV4+8+4HDiBfI4tTm9sLAy/9+HuiMPJVZ/YkUzjMJn18aq
ykerLiSZDJg4ODLrct5qv92Y/LFgeMoPXPVhRGsbBLuIjuHSeZvj4LCVvacoFrKcUjjbiXKuerEI
1u0FTcssuiP1YbKxG2egGgbmThWf2AdO21jGXBPTCvrur8U9hY6KLuFsqTotEQMJMqyqU7U71F0g
LEQTSqqHqpj1SrUVPBl5EPck/9xpfWs9aHyRHfuHwb83Lsh6GstwvFoXMm1rcRC+tUEjGkW/VsKV
fJow8SACRCQ7oCL2m7eNJKPYVUlD/HWaRQ7zeTpcsvnkx9y31SEBrK14DrD4XsAf+IMDKtqmTWPF
2+AGy70nekpIDtHGJbTaS9Eyng5uW1C2sCwJ1coRVKicSuTywJGqdT9CoPAMa1JGOCLmcVnnstCH
hNN2WRPXa3pPJij1Z5GqQxDNN4lIDlx+LDxDmCD9EnG4ZDhu1UVMCVFDWt+kyvmE++fZtuk7WXqt
Qm29+F/jMAQI0LkSx/BfFenFx7xlCK1j06RAEPUvoGZ7WfsyjVPK3HFhB+D9D96fCij0/TfaIMJK
cVjrV/z+11D3rx4Anvd5hH+OuUBFIrrrgYsbST1nmtPP7eKh+++C4kDf0/57hPetzdxtPxyT2Pn5
7vW0DzD7UEuHVsGS2TbVu7gGPlbzZ+yrd3RaEO+BBdycW9xyfQFON0EHLsTl42ZMnBP0uBT9nTPH
lXeqjz45D3+Z9lwbRatah1oDGDAQ0Gq8CnLT6B13pDd+me0VTDWySzcJNriXHGqPl27rSGDHLSZX
IGglSwxhXFxQIofL5VEJahl5+M2nFfwI4uH6ahQU6WUrfbC2akqpI3N1F+t6wub6tmhDpuICvare
5Uo7ItlWU5PA7OO6B/CHgrzPlq+API/FcXVHiBND7KWMQeLTNeOODL7e+ylw2eyXdWKUvPxCr+tA
9C/GgqsX/zDGgJtZux9re9SdVSxLGKpcO8JuMYv/8BVZwMiVdMtdAsXb4rl6wSucHJ2BjPqFatBE
a0d+o9TBZ+SWQqZUgM8poZeCza2OZt4ma3qx+pzJNxIGYrgNRJmQgbJkKB7UYksa/WLNOh1QkzHl
htTBZSH14Pb4ealQYsuVTiyYE0BD7ctGVeczaaBtQuj5i6s/Iukb9DH2oynC4U7XVhHIeZIhRUaf
y71yJ383nLP/Hm6COt1dYnDMCg+duBqp4LCTH5YL0di+r4vbEIzNGQWtoLoCTdbDyDV9p7kyj0E8
047b7v4+YqABVBlAbV7SvoIMkbH8b+fFQiacyMy+uuTfh1tiu0rrRajMCSjeUBhhpzcdlJXV3bTP
DhnoS3DQGpCdeWo7d+egRrqJzHrFogEci2/D0Pq8GIfCBj9SObcNC7DOV8M6Ay3Dt4jvX+bk6UOd
gX/2rAjXSiV+Qs47DJkeT1JnlaYR1gWEcvzOjRUaep71Np3f3Z+e2WYbXpqP4UX6hfTbsU9bJLoO
kHIMWAUSKjwTqFJbBLyN/zTZH1c8kixqeDnkhcpNyjdNRFUY1maUGMuU4kfrF2QNroIbfdTF8k9h
O7DB9mFiCmo9lDkCC65LOJCSE4AF2LrkLCI8OFnMe0VnidzVrphIldE28rgYaHfUIbYVITsBxiEh
hZ8ir17r4uIZEpSRZVJyMJypBTxlxq8LLHF1P+rw03SvXxNYXZNSVF0nE2pU2+AVNAPCBQwk08Dx
0SbrnktVja0kb0ivLX/SdkoYrEf/m99rwUfuwOjkmlQlO+PTUTSa165Ps2E7AHMMwcrAey6nzwuP
Wxu+ArR8+Sa8UA8azgVq0XwfgZS3VmdEvLoIhDKl86/cOEb5XwTZxuIfMm58kyWE71JPj9kTq9Mo
re7kgg+HuCc3QHjfQuk2gobtAnMtNVsF78YCHVdr85phQBgBGMNBrBhNdTDeQYHyfvkcHU7dLpKi
0yq4271AwVU9GYo2vIXcp99cfKUbvHT7/Pv+y5O3l8BMqqg4zJVUWTvwfeqJfNoEBUl0BjY6LbCw
F0pBoiPyhKJat2QM+Cy/A7/y2crct7GEwhkzztw2vKK0nNlDsNbDOF95TEq6FYt4Fa4Xhc1WPZIW
GQdHW1REgGN7qQoDGt/GaJxmFB62pLYJ4ncAP/ZFpkDGb8F88YCmNoM0MKxf4P+kHM/6Pw0YDpd/
iNXmXtyGOGJxCbgJiL/agRUpBtasB31B7ioplHdTsSjKkBzIrod/dAqWL6fy4WHS/fLqVnPd15d5
an/ipTclL4y5KdIOEIBFl9bXxSapE+vTfnkRFpXHqhXMZ4uKalP5Q/YwHHcB9e4anCSeW4FLC/KG
/XDV4rGOwHM7pqaW5XrwoHAAefkFU0BU9+WFSL0N07qW8i//SornGry1wClsm+5EGYt39C3hI5Jg
4r5B8ts7FpHMqT37sL7T3shyVgoe2OCJ/FNsfAM0RZ10ebfL/gsi42CPuxg2cq/nC0U+RlzAMQjM
Fe3OtU16Jr39TGJ9A3790UDE+zsKFAtAaatIgySNBZA+Y5CTM/qQ0XTXNhcsrp5klhhXXeQt5C9x
NXwFKdSGOrzceA0od0RXU6mTdFrxSA9L/Wpp544K+VuVuzEIrylX9tjCjs+LXXp5ibm275jXo+zG
v6R8ec2iwys8Zshx0alo/vKuYluGiPt8KvtPJrmjLkzGNvnNziynq9Vk0LJcFZ7/L0vh6e5hzHeA
ss7Vxuz3g/PyYbpvsY5UuOxXfjDLilo+t+hJfhHFkJWpzDeM2GOd7SwJ5qIiG72XK7KIyZnDw778
XqBnCoWUsj47fMHKnkbPwdcIF/upRnrC3JNRTmn0dghn7MfJOI8sI+L/i82zH7Sn9Xn8cwcvhDT2
mWk3MsjtNyaFI6VIpFE+w/YYwGmHIEWkSNUrv+SAWzIH/3wYWdlpmGCK7wMDgedg2Tv/7R0uJ7c1
45cvzWuJBUKwdHcriwwmsn3Jkh+P9NhzsmkNcbsgrQFjGGl8A8Ga2VAWnlP98Igisi09jmx/JPU3
srNdV8Z0hpxPScGBvX8w/5wS139kIa5Ymx2FqJ8L1fizXTzkrt/khkOi0YVtq3djpCQnx/D5KxEe
Ht4/SloZOsi4nT1fxl9IXTklkvdlKM+K+fwIsSApimk3GhcyF73mehwwZ/s370C9oVeD5Kt1JAI+
vU43Joq7UpnTXI9XUt8vONctXYXNz9R3rDZs2Kk9Z0hJlgeM4nfdex5dSGfcb9o/js9jv5CNWnh6
pfCoFdcr7MR/wSnvuW6WpMW3qZ/hqv+qaDs4t8jtkLuNAv8rxGnLixyYFIrABQAPnFwMAtX0rCb1
7EfwXV0IB9MLxaAsTeX5KVzJSuZr8dBl04rLOJBw2zPTsnvH49AR2xE3xn+HKNzD3e4mTvbu6pUj
89I/eNWyfxrKKiJSjUxSw3/h8p4iOCXZOyWCZ4nPmUMinNVUgkNjeR7xLeoixsY0WcskN0oTJXJc
MPGdBMLl3rlRRCxc8ioMPvWCv8anyhlBS/C233tU1NKa1jJsQrS4ZMgyBBrt8NnmpfQLWM5B6GbU
e73IbUJ8G0G+voOU7vsAn+4F7zJlennUnHrQmuLMG+H+FYX1cgWImr5/uDwWZQBWSmXYdMEu5kmS
zlpfuXFt/kJYojyy02bOyQYN/y9K/luB+txtKiBoYHd8+usVMHBnt9v782G2oec+54fbYUxiFrph
vZqQ8aaI2knkRaVqIIXXX5IeXK3ZzQcSyZw2nrOQsm5yo9J1Mb/CPIQa4h13oWrnKK/JPkAeG0q1
ywL5YXNJaJYPERNHmRSrIYJpfqEGYf+PJyud6xXAG+zcNbUWvwclslUisHBLsEkA0tlukC9fOb5y
iXQABN5yl5wKmFY4oJIiKw/2fuq3viYDJ1sp8j7MYuEGOCdCfSnOxuYO9VDWmV1Uf+jrs9/xMdTh
Q2Qqb7ajJRa2lqORYt9Y+X5NI8CUsGF4jYiWqB4bZeOaRqwf0re8lyWbYD+txwQZpfmZGBrSUvCo
qya9Ftwet5roTQCiZjjMniOVuOiJZLGvDTPvntjrNbToAeAm2+nz3ETShjw/5EPL4JD1N4pjMm3L
UchProt9UcMSSHT2+mEF3o71+r+mgmeBbHqzTFuD5R1+Ey7NZdSVlYxNoLDFnFtlrS72DCEn8szM
oWLt4dZBX34MMXX9ous9b+dT+NR+y2xGW9r1y7Zur+U9nDqOKkUxZomkld7iLnvNxmpN91sOdYAO
Gglc6VoD9u3eHg4POxE/JDu/oA5zE/yY1J61/yetdB3L4Ro9nvonYfs8jf2j9VpyIOwtiaWufEF2
mXWq6dvnjNmkncoKq2vHDphy9MCXhkw+22zS8XADMnGj1GJg24/P+wXdcudBMDLF5YGxCAbQPh9W
nOEC0zw40SlnYE1TSgeIwge1hMk5vsuOqr3i8T6CZE4vXH6XCbO5iZVr9WsmT14F0s1DSvhZgbti
CSqZZeCUv3YI8m+f5gMQwjb16rer1aNKrVqFdoQF0igzfQyMgct9Z4qO+lb/TSV7dj62gsbe4Tm5
Eg+FR4A4iyaikTBzkUdn5qa/jVYk1k933bidB+vwoZvRxZxma+Se3zYAkhZN1p5Ygro/p6Gc9jXs
rKKSBO/1c7RXp6tC8JjjBs4NFoJbNEZEdLnOqPjirRqoVJIjuN2wO4ZgkmKG1rthtBxxhnCYT4w6
YAYSe611jHev4J3xlmDVnzBpScp1sljXLnkja2gKyVdJz7eGDTR4NojH4qAvPLa0fv2biCDy9daq
xD7U2VZNg8wKzopFeF1qF0gRyx0A5y+P1085SxOMZ4CfxprLfs9cN5E3PNNqD/CG0KdNdvfHrbrf
ISkSlYAqUpqn9KlrZM/b/+NXSiN4/NaRrjGwd0a54DVsa2cJ9LP8y83Mk804M4ckHoj9gJkg/cdw
aUv5IMMEmRjgseQa9UGSFslqj6HHBQfriNxDZGsT1co3z3P672K0JBQW8jokxXYAHiq6/iazxoHB
VoKTZ7kw2V58SunTgb2KlLPR5PNBQYhzkgao19bOyjWBdT/2gCVb1HmZa863mXSfn281AaUYtrBm
vdBjdaqp1Ivo+Q0+VLoJ9rwqsW6XZypnVJuKUX/UkYAFO8lZCNtF8FJCjc49q7s1HNhLJm4nA3uW
wsXHgn7XzZlkyNsCurcUKZLTewi4Nv36kagMbZo+SH2T7CpXKIgL+BmJgPb8prbaz3pxE10zSCEx
D4graa2Lbcpn+LmxkuP2lokS3xp+g0Ld5de+dq94dY+KB97w2gZ8yuDwNc7rqXIE47+QKOg92nuc
KAZU2YE/moAFANlZGpdOvQjRbRLXtqthnfIQlzJUjcngdXdXEYw5y+R4HKkn+MQJGJdEcb2nHfbn
qA4xzFug8nlB6hCosAlGU929m5r9tqsue4M9V/GcJSWtfGxalTUZ2kiA0S3xkfT34DGY4VRuhOeE
EM5vu0Qru5C5yGhN1GLThvunHmfEx7qLdOSdGSpmp2HtVm0uC7+5/3j7Z+WjZKJo5G3EV/4JlZHJ
bWLAGPgyjkVr6NM5UCGKut/oXCUnOqAjKtBqQg9Fu03jbTB2gBxJbHE6O4uai+YQhBYlPb1Dz15R
UYLCVIyw8mZa8PACPF3sYu+uxAYCI+qpFnaT0uM7UznPoGO4c0v2eNWDMV68aGFjTrR+738z4ZcZ
sEp/a2/BVSuYDB4MOjtsHhkTSL6iDJiAt8Elj3ptuAAJebY4x6rG8eu4MiL9kvF9x8s+SS0JRewH
8sY6ll1PmjwN1N6ZTOZdI/elGpMEkBvhjViQxfjp3Ks6/ukSPKnHWiISZEGR3AQZypiC696Qet5T
oFeitPpTbIPSs+8G86K7Tgg7+en9XN/o5y6M4dEOXi2X/rtBoOrGn6UWRG9gEttrjyEdEQYu9XFR
4/6qOk3/csqZywpq4Gd+heADdGuc1GYLXFNo2YSkT0EORUV/7IiECk2DL3BTnazKDPVfOe1GyQHq
ib/gXDFVXcAOdNR/FJqZoRiYWZCENeFBl5Nl5mwOsjXCdEwBPhmjsjrod1ql7PAGYYVRtBnZV1xV
4GPeS5J28wUSBd3PulJRDBVSK363ij58n8cIEw6mMwL8EhDywk8Prnqd6NytL05AEnawBLSW6miy
xt13SCuyhOWrsS/hjgcVGvpTOmm3SY3KE1wgtifBKHQMtX3mT4AxgYzrAoiGkPvV0U8/D+lrijtJ
blioxDIRD9X5755bGWbBeVvX6LG05pYKzsZiCWIvdtlvoy8+gzHhrfTHSkBoS9cOQRJBuQqQnHQP
C+tVm9xHSormdlK7eoWpMlmD9Vn0/e9aQ5Ee4npR8CYZPLKaymFu8yKCB3V9T+CIBHGsTVf0JU59
bsa/Ao8J04WZps8rsaGuduFVG31lSpcmJPsLK6uFtVlpouh0JkIwrBCS0UfYScTqauwyiHDvSoIF
AJP5pj3yIgqVvs7hSPfLU10q3yTP2XbYD5nc4PHrADCnbod3jtU7zFVL7zONda/6E3081+TWG18d
Gp42SP3X2w5UiXSQ36U0DgReXjYtLGkuRYZ2ZMZ/AfuzjR4VXirQhdaICVx2QuKO+FjlnrwGmWvU
DhjIaFsziSjPL8QDLvgLmKlUqHnPvFyxsL6zk+3DV1Qby/+uLCiOIaVxgFzHUpXBlUVCLozlvM4X
F37UNeo+/zZA48T+ctFUxH5z/JtZpTebf3tqHoqrtswEhItG61fo1pdZKVucPiuoSnOV6IDQcyw0
N77KvJM5zEx4qlJMcJeSMikErsq4S45wEdcqhlvGkJnI5mE1rht5pW5IXf44byUzsxu6aypqePXf
gc3rv55WSclq+aNhn/Ks6y/YpmOjZ+BVZjvdygAGnD8UBRo35fsHtOazcab3N8l8zEJ9VyzzXdMV
W1n6oPdhx9J35kuKKxeYVM8AywrBgEMmiLf4YVStuf+OUDpxtesokgpqmXA91yHvq1RbE/lXgG1T
NRb7X4/CYtQQVy2KU1HrkfKUEKBm+o8/cqMuhkDxP6EjBOx7mxI0sC6rQ0QFseRV4YhqVctPvUOC
q3YpsFMYc1NIzIrN9jvYSTlJ+USoJ67m4mOZVuWY5gdBBUuLEkHrGdyh2kxLMY85SjFvdwMAwBkR
Qks4WIygZs3Z2zjthSLf3rPJCHlDqh3ikaTu+x7p5vErITdUQfQhK7POKYPfen43isqT/xVufJbs
GCi4OFFqmNqUOjAgRwaOXLPWfr+DUWLVXZkN7U+YkVcIveUC0/xB0SQN+d4rpClcRrFa6+ISC9FW
Id4PSdJQeOFF16oAP2aYbESQhsgbeswyKLfyw/EC82j0Q45fb4ANOoI12ql96Z506ZJ1uG5tz5Bu
fawvTpPiW74mdGQFMGrKuS1mX8mKozp+ayjYv6BlKFq2Y3aOPJ6CZo1qK5rBhtjoFcUCHEor3Yqm
xALAs/1c/eP1mI90YHNDxeyoI7joFsC9xDGgbBT1SnM3KGG2fLnYF25NMUOIVxE02ZWpOfoP0Egj
nPc8kNcP3016Lo8NqfKyG4JOKLhutoliyruEeIxaTmqHTj/IV7eJndkaO1InmsRadV7BQGWlXYqj
jfnonDsoBOKLg7oOQP8ajr0tSnq1VzOFJ6uXnVDB8O5SVsPcUx/zEXMc10ewLPSL8+chbkSQZUBR
1vhf61E3A8QMN0+xGi0jLIaMLbJgWs9X2ZhdzEKAwynvPXw4/WhFqqCQUBbi1PrmP5upNB+zmcf9
LJdZORb6FvCSuUF3Rw3ThWbqkFHuVktJipTz4IQAwX4dz4yI2WHYGSefwRIxA8hhEnqwd6CgQmLB
Ia0aSN6YhJhAdop5wKO7Cdxc4yBdq69uyueC37eF05bVOBiDenGI88RAbDYOd20CHsnLfv2towsE
6Bu8Xm5kmCr8gTPbm5f4Ti3YEIJdphvnC+gr/OrAccXtFhjE35dz/KD6q9aQXR9MYJmSrv8+Uzgs
ZTFEV24C2Fxwd+2GxubiSbphytd6tmTsRpsMNvt1rbUntP8yYl2iV4kTKyikgFHdFjvbwLayNDzN
eFy10RYiPdrzJXv1qwpkj3BxfDp7MLj0zFezdHdKqLd/4s9UtCnvMBWOYRy5HBYMfqF8kwveHX6d
dRlVfllJA4zaQeU9E65kRgagn7EIeeUM20ug+lZrgMWVHYlS0uhTj2NfjCyYFtPgdagNHGrkWMih
dHuWFFL50nvegZzldHTaqAhBTGgxLh+LCdQuyEV3lt8/rNxsIl7Qst/4Ahs3/qYOs8qu1PcTheHE
k0mJy/4SG1tp3GyKfrURWo8kIM66kuBI/TliNZduEb0hx2iTg9vsioLEmAmLqcOanOJd5SRM9qP7
knJubVIYaemm/3Ro24gpZOlCPFK1PZel3mLLHhMmdq/gIvi68DX2xK/gflfoTkcwBPBPMebIh3p2
/DKJvHwx9DsNlzev8clFFNeeiZ7LZNUBZ4HaQbfXxy3iWwd5fnZUfmhmJ/KRX0Q7JpWoDE19AEhT
WB/u+GnnSsZAox/CwBuhXbGlZlp7O0RhhTAuwuAw6PFK+mcfSLEKAjiQ99l+zdEWGJ/gZnd0DiXr
HqMMiwcvP922NcOiOVg8lmATnUYy/INsZO/j6WNN+f/GaC+Bes+FD7aAknG7cWyhZ4wG6M0U0LkW
6pFovOGZ9sgniroopk1qToQCGynzZ8MD8a4c0ehgU5EwkcCjl72bu5257220VJXG45mJDWgLIJji
dQltaJA8RfcliaBEpYkkruRnI6qgz2+MlmYtBoXXVBl95RYzah4VS7RjsnGbCz627SfkvLjc5dDL
HRHXl3wd0Z7q7PHtTeELOqtRzxgNS2PwixX6951ecOTZ0+MOO/qPWUBwu1XS75i/QTe8fUG3UzEJ
gJbDGdMGzEB91AfQMVruCuo8L1cuiVFjmL1zk4xAntxCTRuN2LvwULZQkFH+kmL/eTDY8JR148oj
NF9J4q/ja9i0IVhoEzeSzq1+zdvcYHDXfrQXMVpnpXyPXoVYLpSGeYcp4/LKR02ROQPT/fjKOsa5
fbw7VovV8xGjzQRDkNCUxNSLKTNhS80qPCjNKrZpE4OGOp27WuQ6n9xjpHg+xD4v+TceJQLwwS8F
zyZOIuo+H1Pu8uUobourIjUH9FJMkLJX73FeTVj5owAoB37nRoNPHC6yG2BldgITTXX896GD9ffW
S8WQ4quSekxCQQ8EDHGaRp2SKSRMQsfTp5PvsK90sfpO4W5h3ydJTmqVA2qIfQYAwIYQ0NWlePeY
9NdO1jpdJMnpw7vQANwk0DlV2mdn9wLKoKmqepESR08qzpS81utvO5c/Pi3fgw9lxAHsIvPUUbzt
3QnUyAU/CkCX5QPwNqnxXHdpGfwbDrEzla5aMTbs8XkEq3ELRBkJ6wu/LBivAr9/Cl/DM0SalI1r
ju0yIGtBH6yP77G+1UORiqBOM7miA+TLD1hmCUYATttA2WLvIvUptAg0qIobKwRRhBwf+6a9WW5w
8zerZqvDgPOI/8M0dzJwgSQ55duy3hnpGwOlFTJLcQ++cqFdhEt2Xd0wC61SP8q1CQMIAmrxynm3
VmRu5V7GEXJR/xWiko4wSLGwrVaFdV9B91hOIJcKxU7tPp1o7XKUa7zMK86gHQlJR50ceNWFaiJu
SIArUN6SNKFRlMclWRWYaqKaaj1F2FmTY8JnibBHEUHDH3PCumvAqVuAfKIUmmsg9JPILvcn3kbU
PFi2cLq+1CtELTI4rW5AD/EOPTS+Tr/F582264TevdCGE3OjGcXhZtFdFS0c0xETXq4YrnTRg+Og
wAZkxG+z+XYgAeyR574FEkJrUoAmssnt43kVXFjOCZ1Roh1BhhZSKnHFqwfMlt4B6F+SBhgUs0V3
sTESbcyphUNr1C3xxzq8+391b8S3lFGHa2pXIPNDrQTM4zKZUICBLnL/+SZupSHRbtgyLT00jCn/
p47cxys/ulj1eooZTgPkLbWYd9LRuVyjiLFeoPXmJGmlZP2nuNiSOWZCBaQRttAMZ1oeK6JM8x1h
WGwVCnzMIkWD739z3pdQHD/H/OmM4cUHX9hZC0eNX0HaPiJcOey1AOU/5BFgih+26jF1IPGZmS3R
4h2n30tHse+oopQ8M11Ua8U1QWzR/ffQMF69P/dvnIHZWIELIYgsM80Tw74XJr5AxTKjBzXllxnc
zray8lrHSRRgorUmQnRGSspV22G3S18zJ2t3osXuU0oVNFhdC6YEIOj7gGOYRdpQlvlaWhwOapyb
B5QuEBnb4oN1YIhtyBpAncZOFwavN7DlenVlFtS9M16nvq+R/VXC6/cXxkY6EAHwPv9CmOCNJlW8
PtQ+IULjAF/rERtyKZTdk8CbBHqktowlNxEaHvQpGMxfBsfVSVMXGPRIWkREea4GBzpMAOh0/eEu
xZnK92FLb0YAPvMeR63YhiiIPE5YaWDHbFzQ07nztCkCXTGsBj9T6JN4WXKSp21yPUoeaNOAqwoo
kNRMWULBDCUYn2mq6DqX2O6kp8J6dQ7aLxl2AI5lv0WpnmcvRoU38jOvaQV1WVRj73kVeh9+3D3/
N8FvUv3NH33DnTHk150cHYiGsR8khQrve1kPjL9s6cUbipTUCqHKXcEVf3l/BiKvf6BSgfpfBKPX
BK3eX6xhR5/qMh7WE44IN6NuH5a3IVoH0bo1W9r90zeD3d1T812cpmlCD3aZCTMUZZ+lVwbg6qCe
2b/+967svTJppCP168ApbSckD2WhKdv5M/lehHN6DuUqiRQVqwz1QTtST4XsKCCLd5scAKsZAwGp
jUr40xCONcqAWAt4gaxsN+G72468GOhj1gOpZqfcBd0Uq7Z+y3ZSkDQlxZUpl7Z8kF9GaSoZLarf
XLN9JrkWFffXi1q0sp229itLrswiXLh0/0Mh5E2BGWBHWUYK00qlnezx+AXiVOLhvawLfkfig2N2
gWyBRO/pJPnB9nND/wdtq3fsY1CyVttynBBonmYRv1A/hYDzrJop4JHpOWydf9JMV5suXkJOQBzq
EmwLOsqPwa9HdOzp1rR7DgVKMxNqGU65IAmV+A91XvPvp8MUl7Lt8hFVg45e4dlC/UGSpwgCwipx
PNkdWk3JATENd/cfvREYqXyg3Cadzmsm4RGzAALtPKy95t0Cub4AqCdc5W7M6riibvgDaMHWcxyl
xfiYoc3eqSktsBIpKNO50I6reKhkBxmdSW1WvevoGRVg1RRnrQPUyzi/xVS1d1+1kVl1AoHKeJOj
Prk848jEAeKqk0xG9UIQ6sqJU45gAzeTD6PwNwVf7vnLSh0Gj6oQRCJDkd8+PQiFsawjKCZv+6nf
7ETxpiamE+5AU93THisJttDJMCo9iEHCFR552UHABwqS8yhe7BlTL3PO8oxN1tUKd/5Z5uuIkX34
MLck41P1BOZm1Eg/aHokRClthRRB/4Vnm6qZmYSXpUND4KAQNjBcFjcn9A/TMiS6yPcG7IoZ6Ajc
bcmIdWP/XOwFGYraWBQ9LPwYyTan+FDcJxIQMpOpOvc+6r6zVmUhsij/83zp9ZXaI4QUuMymbHzb
GGdKYsPXuJ3xM2+kHkRWB8t/TUlhMkqVcWAcrsQEXNVCALz1UtG2tvH45V4PacoVvx3owrxdp9h+
Qse4u3um4hdBeCiy5bKtDX4NyxW2DCwfVubOhtAQQCc+QaWlldu9e+SiR8eRMg+BQwW2f3r/sZEK
uyqioqeztUBqH/9UYKbR78SMcuRRsHCdCIc7imZExWAiXPN6bBf0qQBcR99RyTolUn1bOzFMQd43
h+/6IoNNedinCrcEdTbEJXQUcLuIgcUC7YEzOhGvDNJeK0ZxBE/dhVmY9EMVMxGu+QXnwAVktQMA
ulmZvuJshe61tfmIOAYjLVjyxhrtjQ3J7gkiwCGPhsAuZ9xMdVbSd7je5Br/6c3ILFgF2WkLcyZl
UtAiD3/UilAZ890aS9lvFUqPfYWr0BMtaFotWjkoWL8vyKfUqyLra59ZG+eUIfKG8epWXJ462R8L
RCgRMlVCV65TRBMAd45M52GdkfkSCLX9Nqqak3afrpt7r7EXAcHzNh29HphfCXOnJxh+SbRzJsUY
UTzQ+fOoueShy6jrAIHVw368xY9gT72mND6jsU8eCXyn+8iua6ynorejimvLM8yXNAnFHkNOdNrh
PrP2CVjk2Ohn3zWHAN9ZGunrLRENZijljcMX1Ee0HQz+s+C8Pw4ksEYQJ8QEp1KEAGVlbBkC1o4j
PDSuHX7QTduoCIPh+wWDnb6LOL+QIGsEU9NPyZfa+nAu9TWKXEvlQKHmzHHX0Goaboe0awiEnK7K
jrcFJxp87uk2yiijbb/Wa03CEAbnW9JTcrY734wRkiwQVmZj2wcuy+kHJ4XlOaxoBCIvU0BlPpq9
kU1aQuIVkIfBYqxpT2Df9Z3/u2mPIXB1i8wWso3W2BQyopx65sUxsw8fyMVVkDaBrQPfA75zjMDF
uEcwK49acent+EDAtGjxNbzjILG5LPXITw9WVx1Po6me20VdSGv8Yhkb+3Vd/s4s2u0P7+Y4VAp1
2v3SOWpvXejoAYskq93f0DiyL4xnL48JVBhGHS74
`protect end_protected
