-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
eGKIIIrkzhjMyJq+8beXhxbNj0KyWRd+ExAUpRmFVq7WIj9h7PjF0Z4QIPau/WFbcr5J4rNShkg9
WUUXWDWwZLaYZF9YQSiCVMYuHcAtIUoBwrTTm+tnvobuX0RcULv30OrQJEYpUM+exPPUrlgTnxyi
wHK//gzSIN8a3PVMYEm1AFDfUMkJkrnJKKDXdd11Oz8iAqpk3nwdmNcY+eP5xyQUhmI8J67Cl/iM
4rVP3k/tn7lwGZjH0WhiAKxMot5KLMlnhCdajwDfIZUvpUqWjbdtoJI+ZUCjj0ZoaqWBxN8SuB2t
0+VTT044tngMx1zqorkWGeNzKl/W1X4NvCrMTw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6512)
`protect data_block
QFHRqprXsBooQqX4OgWaPPyfvbpuqoybNL6qX9Njd0Kx2kKHOjS69NRyq7lHh9Kf+87rvnNrVQTH
3Qcx2romKHjCWc/v4V8iBSL/Tj17b909AQToJhPLW08GOBl3lI6GKWk+I9X+2lxaDzlNs6stxVQH
ITBJzR6svqlzDyBZr1z4tYWzl7KnU/1OU01x+oldjxxBpICsTp7PZmaIrgXiaMmoowmQ52ur24MI
9qJYpVzroQvSWUCpOxRC1wC1CkKmifvXa4+O31QtVq79xxFNZZSJ6iYfEnCxfhSonkBVG9DROfuZ
RUkbNiJ7zk0D+f+TuQiYuWcG2lHLGcf8QEztYdkrCfFIJy+sM+qnOkRR412etl7Cs6lOvIPL6WZt
FJQp4iY2owL4Qk2gzFQR25ZyzygaRr4Jm14/spyPF0vET5dplmbEzNTgPuTPUlPlzJdliZC4BM0q
aJNFbviLv3OXZ/IF3dnEVn2gSyYdX3IbSXXJXfqMdY3AicLo77SCKXlW5+xJjYLd5HJHoGp83Yl0
ydohzeOYcHwUnzVbwhp3oGZYKqt3w5ihwYmIfiIYW8dsYvLEjZXKZdpPVW6XQBbobCblncOKxyqD
TvPincohGJ5exSKpubN8BH/7B7NK3UIP7nr1Be+1x3crBMQrQP7ltjKAoHiRxkhjq2hrV5v17IkU
d9iRSpdZW+yHi+7q0Gs8w1EKIEs+WLgl3JGJ7dqE743Yx//xV4QQBuF9eletxZW3myN2o+iujs5Z
ZtXqVMGF34h8DSOOydu4UiWRmCKM3WTO1KTlxSS6EJb9oujdQczvmWtrBtEo75VvaQL6W+axGeld
9nWpfQHGOta+Bi/9QcodFeATKbxtvd0Gvan+c2TPAfAT563irqsot5YeeC3SXrEfVcoLYqvcr/jW
oTkpH3uPwN36KhPtXL70im/hXa2q1Q0LX3EiaqfhcdneHSiEAyAe1/3ve37B2bXkDBsx5Tj2mo//
eLYAD9rnoiE7meP2L6RnkajFrJqCsNVxhXjuHoK6OM8Fuio62IEb5674lxZseAA74Ntk2qIYR0jD
gI3Ml3S382veO5LRjU4W488dNO/Yd2gRRKJ8Hp1qv7V+GDKfD5AwbVdxwiPTiKUaiTZHKyB/tXzU
dwyyLlMJ7cwKcWmq8bmCHXEfyer9BrOb3QZANu3aF2zy5e2P2Ewr+C+v7Ojf1neojklTl08VydqK
vf8glnPPj0Kyild9hRp4rgpl81isewmAQCiNlYbNHGv3/YNIlPmrcr93kCaC2N6Pk72JlNq3g7UX
xEcUBY2eEaZlFgjOJJlE0eLyILSPImILF1G06GdgS96IR3NhomR8ZT9zBM4FWad5i+FczX3R/5Wa
KBKe3tFoYsakIt61HRMPQyNL1p787CYRJIT/vGde8hKJVNrQUCezCmDHrMhKBD3UuNYurZjpcue0
Nucd9LQct01RRIRAs+Q5ArhadvMJqEGE5mDrndB2Silvc/bfYm1y7L0O/IgwCeyZnGlODheqnGSO
Pp5+A5TKVZGMGnV89BRhfY+QWlbateuNTD7JRUNQv3ilhRxhvMDXu9VffH26n5hQnC8M1Ds2H0yq
jclHYAIPqYlwrLZmGxGs8Iqk2owz/4gren2BwSO3wmDkTv7n2fxnKTYiFQFUwGQVWm+gN7FpBaHs
mLMH9CJuWWybHFU2eh/YlmgcjJDc1M5JWk+tp5ASVnRNN3JSpJ8KoSEP6mnbjVe19erJNvfxTZWk
gghsR9atiswrW4xHc9UQJdVm9bEQ5TN5PnmJe08PI1s5FLqeiICOVYsRo86FS3ojM029+hCo1JFK
CWfwU454eOKs53539AdyeYKYP/RNaWE/1NhJZ9oB13PVPG530YUd22841mux7hzfNsvGs+fKCTy5
PQnw4uOh9/xPB4u60HqhFgegeQPI7CotjVAC2yK/t1PvQj+P7Ca8det2Z2rBtcLwzWh4zQQ0QHVZ
rERels443irIr6S1UNxNrJVfNpmSJOLyNZhVb2CpWNnbFcDDh2NSMSF5Gak/Jy/NviCo0VSEhkE7
7NUcdYitApee9LD5l0cWdB7784KFG5YEAjf8VBIHtkMuX4O8AqYI1XzdbOC/zTm3JAYkgxL5z9mM
T15GaNUUPveHojUNVIHDR/oFhaQJ4yAyHgmiFIcY7/HgmOO74VqwehzWDK5g2zT0yhhPX9nI4UsE
g7hjHTNV+ZqfllsC+e+r0HbRflySNk+c3DNanthZGZGKk9XkRjBnr2H71hD396IJR2LFwYpJZXmu
hH5R2mtt1Vr4oAsEsPVXUvcw0zf3DCuqZdQcwlBJxBzyrr2Ob+hs2/bM3b/ZU0k6/x8yZ1OWD321
8yHmLV+0aA5uglVzx+lWn9xDICMs0lUnNF/lzATSrgt/qg6aQxbJ5ZrCh1KCaFJuXaSSAiaVuMHH
OaFXFm9NqBHHWHqJigJeZ1Oi5sNqpEc1Wj1+xS5TSuvGm+AHJ7nBlkA/YKta1gOrPJ1WukuKVSFq
9EdZe3LSgmE3cCohwX3F43VLXJdr1Tcct3Ksep0RtdrcBI4H5cQrvE4yG13MnIPYh8zj7UmjEm3m
0lFN6lHmbrBYH3umCnKk8aRJmZvz3PQk2ci09onnBrr4oVkZkVSll8vZGm+SCizmUTtj1QdHq6To
LYegr/BAfkF1OhXL8fyXcxjuacwDmJkXpmphr/Vz9h/DypbXio4QJMZW0r5wKzrOEWCWFSoxo9hw
f1swl+jiVVlPk8hMY5VlyhQuaa3GY9zNxBq9rgTyaeGpXVoEZlI3J8qinVr9CEI31TKMpD385Wtg
gSYvLXyEyuyDN1NSvnDryq0BoBcxvrNA4ObFK3KRIQoSLZXvLoOVjmhBRfNxxweuqGJQoBTyjbkM
wy1uzFJJbFWoX/BcV9pQXxe9HacPpr1laf965VUrUnq1JHnvANxKd+PTdlaLMZraDwtydtBwTS7E
CM/pXRBLogQd9jGPf/y1IMaE3d38tXcec2AL/fp9mF4q2aUUoSdh/LRmGitY2wEoISFly2U8iDo+
4GEISSIaV+eZoxv7M+tMpPJdHCa8tUB/jNRHOBDm+780YdKd4ZEQA5QUthW5+WBrzBSpAuz/8Zgw
ZCswTAnCPLc9IQKt7ghWbXc8mS5L5T9HMm3x3UiM7hO4bP99DzsCGtMCfjNcdqGgQAEQGQV8YpiR
i0VcFK9Mc5pyaUxNpalJco/UQz4fTRuMxcildfUfgwmpt/4DHIBCZVsNwwLfE6NTbj3vnC+0IOum
7mpIfg0E9A4VSMBkf7FyBKNUv6ezKpuPb47SVnvz4aIyGBku4ePd7vGIev/39EUyKaY/rWwjqccG
ifALZREZHA809nN9FCEjm+I906apW0WMjdBqVrvliTGSgDrWCwd0nZZMoxRRGs7wi5AetCG5EVlJ
M6Do5cbmzISvoq2G+RHXhi7scNYftdUcCDQjrzLeU0jA2Iow2X8FNkR54eviCquai4w9Z6iTBP8P
iNqe0pT+O89IxQOgsdm4DwAgzHRgYbXT4H44sMmwFYZNLh3+fXPzBkuyAoq3XJHXuDrWI9wrh7Dk
RRVoWpwc7kPoda7cAJtkP7vtXjDlHYheWAAVVNoDwx0VrAUcy4TRbaSVwGz2pyMK6Cno6bB9INJk
yXVO+W5xvtFO04GmiyXK5PERJxyvmGJk1bw2mx7C1sM9cAIHT7Az5bK2GshULaaFHb/YsjHrEWqF
Y1oIrCPCXE6iD8lVm+yfzUDQv23qv0vyqaRY7iJ4nrbD4WXTJZF2N62ZliJO6Wsl3O3V7a8ie9FL
vp33MzquLhuVLOE5tO+YJ4p4nVTVDWcx0yXimq6DBF1pety0NXjNuTkgFh8ngztxucnq63lMsh52
fLwpJvf6X5rDvQbOZxeClmptFRCp9Xsf8tgUcMQY8t8FPysgs/096oOZC2D1N7Jk97dFph097rjl
AFZjK1cgL8UeeE0pxf4lNbIqYS+ZrHh8XaFE/uCSbvi+k+B8E1VTgnz/HnbKVdI/roZ1i9E/2RCK
jmmyHoIIldzOnzFrKNnu7UV4FGUjdAD2AaRSJonf+yscdzxW0poZjMpKOWtwQoRWh+7lg0ytGL3f
5T4sSnhiWy3+jiep4bABnujbzCbMyOK/EKQtc9gi4GLe6igZVt/VzfP7vNA+xgPNB0gBZwPa/Ltr
6L1zksXWGf2bd5Vk05I2pLKZFsepuiVPvKyEPWwhbKh4wMKF8Iwm+4HUrB02E/eIobK2yfB8IlyW
ut4u3+Jklv5CGDA+cYY45crmetcWBHmV4I0I7rSVLu8haIHih6GSlvVToqw8/qHpjhpoLepaZli+
0y8fDFF41Uvqx/xS9hYEWu3fx0erp8dJHD9dQQDrDEnJ9fb739XD+/x5rh+qle++lFizl8yAt69A
+ar02fIpfLM+DpLtDG6gAzxUBLrd+EtXPZUMmKREu5kHrWovrgQ0hN+2TX7Zao++nLh63IkoxoEa
oOw6n79aR4P2MdrvNeAEvSztVJ5gjhqb3Ipi61HBcjjrwINWfVlCEWXfHo+f6XJ/Y8RSVyoI5VIE
TOaIrNGlCSuRU3V/7CBR+740UpfEodA8A3nP/eKJhZPOfP8V2oi/i7tD6/HzmUTbbH9+hs5RE6QX
eppn73xXzr+P6pWSGDcNsBSbiJv6e4afE2TmjKdn3N7zBtvRLXiw8pVNq4f7Z2OLZZC0a/0Uh9U/
kyoOi96tyqvweM182EUgoN5fLesQKukhBuaKy9N8vl3BtuPPh/THIKo4jbkgEa90aaJNN6L7EW1R
wZpO70bt0fgDbwy4S+B5fGRmiI1jG4TOl0Ezz2oqG/IUNSlQrIP/5WSfDKFzrhv8wV7ca/4JN/nw
xhvhmthsnlw5sNTd+GTo9L4FpWMYu0zSKd+5VhRCI0Fk/yvaSzBrvvSjgTcPk14DWuFEFYcj13tM
QjzXvLKTcDSYQ0qAbhGmjSWiHQrwGVXw7FdbYzWD715iwXtUm+knG/zFkwegMpC1H5Pqn9oDmtkX
lEVfgbu2EcIoCiOv6YdFypfbEBT5RnfDcJ6o2KfaES0xI/HtwC9rSV4e337033j9w0pugPNTc0dg
nTY/Mr15wkV2CaB2p7bJSLPkpIUY4OsvjPks2i2+FZfm7vUnT9z/iz2f7KwdkKM9WoxRZFicaVZ8
iRyciEtp6ERdb1XFTt2pVvg3Ek0mVvNngMHQcz36Xjedl+cbJ1dB3dejhyub73RmQ7ZwYiltH6qP
x/Df4uDV83r23YuRE11/hv7hyDBFhNf9M1AiKh1H3jVvXT8SthHURns3eNAs4G+cn0f2iS4EF/vW
DEyRvhvMKR3q4QWco/EnzEPCawMfvPavlOB8pZW6YTQ4+BFqK6zF8TFFyYk5ip77+L4LiVTqKPMc
1l8RIbivAxEQ8Oyo3BxWebBxeJNEFSZd34IZW/YGYUD4kM2a6zP2UwPuHgCROIl1C1X0VYav9Aiy
OGGjIqILccF5OevCzwTtI+PFhKm+I0IELrVeVGqDIlv01RxZp25pbFB7mvkNOljr2JFVKGJ0CE0D
5KvoWaImZAaTVqYWp9kBNXX2k77Udf06lfK+M+dzJw7cdtRJ9xV4Y7twKvLUVQlAqXLGH80PMoFK
IQB8fAhvmXUSdrxAjIFJ6bWYgKgL9JME8PHHnyd00UXJK+4lZIsa0BFpWuYTQ6Ht/svZXJjJp+lj
CaL5N/wBj72lLtjKPwrbOS705YBk2tFrbcp8S1Xem/xPs+UxbY/Tz98WkJTsP62z1tyZVkkQRh1H
Z+OG0dMmlFykL2L4N46f4ys9MKAVkUXclwg/gwMQst2nRMy9DRvcGKUfir8OkyBYjXZ/jUSHZZX3
cHy6EkQOGXr/6aTfxUkk69BBody7Nym4emb48io73M9iy3zp6fuFZDcBYqLr0v9W59vaGKfeUB5n
dfmh2e/9QlNvvjPppyRa5jA26tVpJVeaaJUskl+1kf5Aq3ENvovJMpVbR+Kb/Ukom2pwZK5uTQD4
nFkiaz22sVoPJo2SOApO4sV256Tl4mcnmKaLsQDPpfU3qUTuVpM4Uw8pKHk0Bsv87kT+qFIoZQ4M
olwsj1oOcWBKck8iXbtmfHdBFP0PxGeV51SqL4Ekm3BhPmeFp+ALyzYgap052wZQlu8kHc866y1L
zcwJoeEHBjaNUAwVAkSChoEAgHflLTubn/hujuO2w31Sel1fqZyntv4WVaMMalyKMabTpnW0LkWD
wxsklqTv0GKk1Hv8wz8GqqshokSNqF3LrOMdt2poDpfazG5dbPuA+w/w36Xk8oclFxaBNq53BvhY
W/0X0kiiBO2CnYJtozHneWLToVUiEHKBJSG0DcIetk4gqFtdsQ9xuJHbbISk0OEfItUvQWwnQxCj
5Iah3Bc2UtAhLm2jwu1tCMDNlgpkDKv2p8WczR5U7+QKaHykR4qwKzY0bcw+gpOfYYylGHJumnjz
r/T4mG8Y90eXDX8FqlAW9eXAsiDChscyRyU5j7CsCqLUnMwprm4SRYQy97HPSGivQvcDn0Wzy6zt
v+YOcz3Y8BmrbW6Nsvj+DRlAr8Tkt65OGd04nSH1cg1DuWGTR9V0aS4Dxd8OYfl5CORgAKnXk+Hw
jzJz/iUUIYPelpBpdA4ck/71c2vtyZ/NS+DzQsWOBX1f+TdW5WcCkJ9/vX3BHU0IyV3NJ71UbpBN
gkX4gnLoN1yrHAeeCXrkzWYtTwTWgjrBdUABtDbe75kiahguEIJ8p0sJpFRPr8+3mxsxwozWdcKX
Wt4vdOsRg7ZZbWrGe79hK4lG7mssDs21gMlpONDLna5ZHUYD+ZcGu2P/G5KhobMdopzNCrlLuRO6
hx0jSB6tq8m4wFNa4x85pDzfv2uAf0NwccwIfh+29K/Rf7m0P4zeGkRmWIs0Ybi4wUUnp5y4jciO
Ee+sYZU4c84JyMkdgAdUNGlx0BO+Fb5nUsGzkZgBpeGUSb8QDaRaPgjhD8aPhIQCpjt5o+zPtLlw
EujcxNL4XCvI3M2mHvS58pYiYcPjgWNW5muKCOaG8TXswH53ojWbbsUJCgtQ80efVMiMcno30zjF
c9eMan6sqH7Rkq88Mwz8layIGFqsr8cIb/4atY7npCwzJd4y+SOde+FrXgcP3ngimzCUe1HWWQJl
lF8VpfqBomEJh6gN4VRygrSdH8WZqNUw2hvHt7FFW5IsUPKghRFh3h+7mUI/2GwQtdsieD4AHiJm
IlL+zZ5mXqnaqq6qnifGBsB3mAU11optMk0u/ZhfqWAncMeK734AEwf90cgpnckLq3X2cRbUK6zV
yLh2hD1dLr4Fx2EMop0qa7v2fsjQE3eYXOZCgRqQRjfQ+976n470mW4rcXHzGUisquLJ3WAf9SdX
DMYlQXIBWDf71Mkcs7L9WuhtaKB0SIpCia5FLHiLxLKCTkmVt2xaDzJ2RTIesINYJ5NsrXW5eqRY
dsaTqP+QRn+8XhzA0ikuj+1d3WJRXHJ7ZzDBkS/p0GIBvk5CQfAvUhVdakBrCAUsc2PbR+NQGq9G
IMdvVfXxjOYnjHnUIv/lH9h0ERwPTWb9tK7cG6zsWnDzFvb7bTTm0awHpEzcAd6Lk1OYwZz0SRSW
2VwQpWe5M+NUT2jYzq02zAcKtnYf1ManI9sEsdOqmkm2iqBwJeWpKbCELk60lRkepftiyfXAAtM9
HjqaeaoOnXm+/EFqi5uV22WrRXqyQruY+9k3bWaxVAsq0FrgtTi7rmxNlgKXr3HID3UGFoCot6uu
HKMswV3BDig+GaaZxTtXtC1LRehqj/R+JrwA8Nt0Jq/f6h4x+68iQvgzznp+cuS/Uq6lhkA1URWm
4/iHJ4bvV13OsHA6o4B3RjpTmR/7zVTRWSTHsruWcjTRloDHNuwll7HVThKiEX1cLVSAQxdKrhXm
XLcBNdXTT0+eYAtIJB6dZ0uTPOGoRV2VdCzSKDApq84+B9Gn3n1IrXo8KijKo87PWJNwlMtL7XxA
IOR8tFQLtt5OZoSryxRZUr9cF+CqjY+rhgOfXABAdouhaV4Wq98UwyDR4NMufCuAVThZcY+z/n3j
GODhH0Y7N2GBCRwPiPxo7Uv3XstA/T0Q+k/RXBaLavmuaX81Dwq1zKbmcoQodE3wEwNUdxslVSHb
L+eQ0DlQ2BXM6QRPd/rtqrK76e6w1PldK1qaIUPvnA3eIl7uca7zcGUsTZpVHktBnmZ41N/gnFTQ
jhvvcoIaqjaZUOE7XTiRCYPfXoEMzZl3U2GizDQB/9KEVHPVKQjoGEKx+vn7afEoe4jiIbw6+K30
d+1xSXYdnm88eNXy7COR0yc6XOdXdo8qAwEwvwsx08pYaQHZqCXpXZIZ5RsToAhgiuc8+CHbD0pN
cEeWF+/xJ2XKoNTzHx7MeQWuiE3Co+23AFOlylCYXo7vtWjzFcsa+WqNCy4zrykzrPv7ncm712/X
1if856xeVqJfYWE2O32TeUGa63/TmoWlbwFPb3/Gi4V5MZuLY5rfY6B6Yw92UysIOo/QEtOE/YUU
gi88B80oBpvYg7cc+uXsQmcGkNAfYwxkpOUy36EZkc42srsAE8b5Gesa1WCSAdY1Vm36zYB+SpTi
Fynflp7E+Q4LloCUNULwCFQKNJa/YEw3WveQ0De5HMMAgWEaDVQ34xRKfsGWA11WLVU9WnwkIB1i
vD0svKRTZW11hD9we60=
`protect end_protected
