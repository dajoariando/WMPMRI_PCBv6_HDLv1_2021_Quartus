-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
LpjcFmjwz+8/yMRHrAi5jLaRzwHSe073MnHkcaJplo8fpYTm4GOXQ4tfPlSroHbbYNXokVLZANgM
D1JBAGtGyhF8mUMVV9w+WxQxVgG5Ah9OeQheROAMP1XYM4pb0ZT4g3a0lfP0xR8S2eRl7QnnVvTR
cr/9wCTjtIKeJVL1uuPi/O/PEfRD63oHtMJ6pVDQYCG/WIwTHFiIkrEJU526+Ve3D+yBzAiW5C6B
dSmhTGxbSnijeqsgE1Efg0B5Add3KyIBQMhezkcrHKXHf9y52WIA4IZcZAXgqJY/O/LDJquz0SFY
WNybsj7irGUg7uW72LYk5A/Omt24QrFUU2Ryqg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4288)
`protect data_block
CRqW8Y34nSfSuo9Kpqxt+vDYQshbgcTxKr5QnWCJQa3C1E+VMM0Vtw9UsfepDU6GtgLyB6H4S9XM
dOgHaHg/OCejttOfmcx0s7KizOO3UEXBTDf4PPTE5VD2Upw6EvIkquJ2EsuIKMIRczQS5aEmCBIN
eM/FCKizQ5nr748klm6Vf4dRM93BD1Lfzm4CZtMcL2L9+wN88cttu+/90m6pGwAZC6KxdEVUzklA
oA5zF5vprqzcRHyLjdyz+AVOe46uJ5MWxMm2qUulJ068feO2xjBOk80mSgzDr0yOm94JhUoGP9Ix
S3DEIykkMxTaW/RoTBpeIOsxwICY2mFTGUNLmASTz3F3fY/zggNlVPv2b0oFbNOwavM3FNJ5Wxkc
2nqq0MLFIUe2XV2TCQFLjUP/mScJhq+vqLikW92DTFjz/jtYKysA9hD4lhrg3M1V69vD/i+9h2Fy
K3qAFJ1xKTiK3wj3Ne4OzHqljM9G7gXzGC7KYxsPWO3uNBFIWfVuUz5JWFi8loSkNlgBUVYDhUMi
AhV4uR7tbRvhIBYrBNuireVEqj4bBgETh3jvslJm/Z2WfOEa+MwKaLNeCRwLMfwHR3CLI0yxM8S5
JcYOoePAhr9PkusXdlVXXefKLUnqykPxA4fhwXr4+PL256qRsjGxrCUkM/bmjnoFF6+4wxsHz6Tw
IBCL/Z1g18Pevr65JpPU8KoA8X4k6fbNPXJh2gfYeTPI94keS0F7Vu6oeHO95Jp3oV90U7Rn7Y2a
3ZXizt5xYUJa1kJttb8daNj3dudDQcGga3JWEExvOE7lMjm7RuK+Iek9rg66ID0xAZh6YsRHTyMN
vdTBcuYf0vo6TGvdxLoCytkOdCu1XNaFMl8ScK7SZf3Xnbmxv5dF6XfRidttsvjOJ7eTJaVPibdo
BuEVJY9J04fpTzOQyZIc9xTSBvJiqfoxcXfSGDyzfMfS5Xkn+9XW76dCsSZ/ooumKUPIislypLNR
FcU/0Wvmdx3dBtsl85JKfTroyk8D195c0RBLYSP3+VOdz+gxDiipZc6wE7wi6uguNrpWcRoz8OFg
17pQtiMh6NuSm5fAYk1AYMpYQcEIkEAwOJZFMQ/bdSu98ntsJYu4bSyB2yNK5fG3+QAsI6BYaBdl
qRl1e9bkwvjb+i/T/W5Kmp/qSycOeyqgT9Ui/pXWapFezx9pAAzMzOtEnBvS7PGsz/iccxvIKTDt
TsxMVJC3LhFwmmqJq/4r4BTJODq/mI3uiTP6/ivCJigMgZ65AwyDAO5Xh6aGGaHSLYzlJvkipvIi
GeUcqhOLRTrx0GhfF/WpL9WtwoQY3qB3V0va6HhgumvVRbA7VfwHdfNm1u1zIf0A8FvkHobrYaMG
acZ1O1v0jhmS1rpvnqwHneGvLWTvlSwrE80/JNLnUqCZ1NYE8NIDQiBzrnsErnqkqei5qzj5Cd03
S5g2RUFC22Tph7qoizZKEw0+4+RT/iVbJWKHXZpIJ3mZmIG5vYviAqPAiJuBn0G20aMBjXT8Eaau
U19KXBL7JfudNyHaCz6V8IOWBpc/EDc9+PiaC9nHv99Q6+DCBcEfwiuoLyyAh2mn7/ANsAoeRwTF
ONnMbreqvMPvzeidug3kLZ79GJ7Itpug1Lk1iDIqFPnMQWy0erz9rNXXvY35vZ5cV5aGARa0hTJt
7a1gmCzjjQQ2IFiqtDoTF3dq081cebqpD5+FTZ0YCDsFlxiVNufmS6itOws+T7F/eUIBl/gSCRee
uNGgZZHI1pfyunrVk8Q26bS/SCRicg/QgY61YTL5csRJpS1JPtBKHNwUQATLHDfGx9bS/asRDYoE
OeI4zy/DKIDsfreZNU4J4jwLheqOEvFCl7UeUnqrA05+5Kj7fqIJrTYyRnYB07lkhdNM9kdIAEMY
Z3b8e6mUwH3E4mQkMk189TpmI3o7RnRqcpHquvPaKpA5k74YBT/iO0pJJ5dlkBSG7jf+9kZtIcmb
BYOYkRpIXzA1nc8J5TTO/7TayvlfWFOg5A0PN2/EWfsQORkVJ8ca+Nfrx8E0w3eS8YmguNXUroMa
At1U+bVeDkHWJVD30VSpkZ0r7kX+4uF0jNduOjgCcyUwDlCMY4XnMPLJBJn9cD61HGvETMZhtUXg
7QpPcuk3gReORlDlTKOZtkQqo2q+mEkPOzEjB62qBVO9taRwyLA8Lj3x10SzoCJ4XvJiv+MBuv1w
9/gOdnDRdFh4HkkKyIXWx7BRlp6berqurNpcId8Lg8icVMBx6FQUQRa0JF8GL0S8rgswyBAOCCRG
4lFRuJIPB7FLG2ZMHufnbKq5oVNv7Mt8aY7jtuu/bSyMCaN+9cnRKaRDPtyHw7RgGMnVeFAb0Vc4
Nxe+UW785isacxZ5naKbVz3ngfUP149Mt5QN5E150ZkvXq53DhlXZhgDjyrZejPH4xkkd0mSiG/U
HmDHQ1F3Yi67IEzJNFngvAMaJ5EV262nxNYrRsw9W/IQ1GqFVJ6a/zv0yJzd643N0nPy4Tl/I7AY
DRzCVdhVQRfK+wde1QRswNfNkWLgLAxWNHo8U4EtD5+ByxTJidZN9h27ZAiOPwc3Sf6rE/iWs13r
N9EQBrPjKrEK3+EtO/R89/GX8s1nVNJTV9J72wAqv7YUOlRl4HzEK9whTKKYkSHrsp+p4lRhN8pn
kEHkxb/9dbkd+yGUZvXRhErvM4Sk3FUIqqlYnTPe7QF01vmjeTcpKT+CpQ6Sx6oe4vyIY+FHQrUv
vcGJuhgvlmWaeV32HkgraaA3CpE1SmrL3/rdyA7SlYbjxYWH70mykS/FqMJChBNehu0+jr67ES1D
CClc4shFQVEqncj6EqNqMrdMVw3Dh0n0euW0IAis6iQ3hQIYopBwlNUYqX5mUvYvQ6GRDTrg8jzO
AGPKvuM0bNTNBndI08JTx/s2sfTebhv3+zkU4prQpzkiFGN48elhtifNEqS4x2yILIJXTvuhELxg
GyAqm2M/VIdxMyWhqMJgtMOx7B5tE/MY93y5EKZu0JFSISkQVJnO71pH0CIB5OO8IcHgP0UBl2Qj
D3drdaZ58XR75DnfVd5oMVJJA5mHGrpQ3wMZ+o613xXSY+2PO/F+s7tN47lpvVVVIbS/qrUqmRph
I/FJ4IXQmdrLWKkf7vpgGhiRUUZ/H7RIXTakRX+9Hlt0g7rAl6+zC3hYMK3ceZO9CSgF1R4Wu8Vh
ajhhdkJ8DFc4BN+oWx5xviGqSYXSbL/XjFPZX/RS+N5TTyMRP6FLnXDwY967sWzb1AD4Hlh2PGiB
a5NrN5hkLz27UwY8WdhpS/05z6XiIre2zCkNEaH75z+FbMLEzieDJC29f/vIG8a245RG3FB2+t7C
z+DYDmk4Wtr2PuSs3Qk4EIAFgcvb+cwDFmV7IE3GPYei82KYDIkd3YmK/tMtUwwbZgYKVFkMWDXe
5bkldrLve6B0vPrrI3o+Gsz13Jt1ZhBlIpm2VbzB8TK/o8mD2wivys9v9hTdHcBhl214gkTY02ak
tsKrLX0CpKMb6FpgVmVfhvwTuFGlriG0SvZI7MbouU3GLRE/STbu6wNuIkdx8OrlCrLqacE5qSrr
LI46DnSFB6wY1LimqNNjAk0ZMKNCvpckCWDq9Gw4jJDKnru9WXhOAjl8CbFPX+R8qzW+jIWbilds
NBErX1p7BO58MssIktaiN7TAO5aHwXa0UHhc9TFjCr26UXj5VGU4aZwxeBZkXMmbxxzWQN/4R9aw
VJBm6+Q3eZ00tiZloMnyM01Hd1kHuX9ROZ5Q1zrHWJg0uQNfGBt5VplKkEKShSaqqkJw6BkFH3BK
PmSc3SypgEn1dQ81pD+WARD+Cby3J9yp9QTLo5fFWSc4chkmQnq6VJPEiAm4UNEYnCXmRkwIFzG/
TNAiM1ubOuuahnKtg+z4OipJ3PMZ/lDhLIm//y7J+JsSSdKhaSJGd0ai85J6NCY2ip9U40Zvlg6v
90iSpVrTnrKIOx/JdDNbZ02LiEfwhKW6nudn55Y+lhK4KMJk2HS1K3BUegum1e0DIyEUKVgSAB4a
LTC32QfExgwUrpFG6XYvrhddoKRgSIcOfqXhM7dxZD/DR5A7lWApKQyh1ybrbqwmUulsqVEGa2x6
IIapZjzh3Y+nHnrZxJQR4z96KR3qUhcx041sBpAN5WGdaPkPXXG7/cqaKoUhzg6ecCfqsYNYxqfR
kArKNVZzLntj+TEq38Sr6cuNt4XDiJovNuseByBO2AIVr9+FDidkDmhI0RgYFjPwP87bCmAgTgnl
sNazJmU0TG5Bway9+8mSwgZDgsItuoDIGe+5NlAqGso8H71c8XDyWI7+f6inj7yaWFSY8ZYZDnft
H4QiZXWyO/fvY9YnQ+FNWFv8pDbA7RudP/gupvV+L/zMxvb+LlD/eE5SV69g++6k9/bJzeSU2UV/
vzxsrR1/Eah1M5V9IKwTFYn+cHAaTHdYyC5S7C9ovL/7vvAO99P/Wn8/oFIinitpcuRVWeAU9gPv
00+BgKLZ8PwPmOdYpFMUVqjq/QvuKxTtpuBqqF9D3Ps3zx+qJJVbLTzx/N4ZkBwqbukiq35QgokH
SIPrkd5pfCtRKmkO5q/M/IOjjhZ8O/7laXSyFcUQeOv01hlEVIGfeyHP6Z9cLDjhCaJAE2gO0B8k
m3pRN4yJsRB3fwPt6rYEgewcjGEG1l+wwF88hBCAJ1Bf8gVzVSF8exYztXx0jHCHJBTj+85RemA6
A8vQkqrqluV3O1w72iZSHiHRwVGxiWPxel+WFAVH619ERMOdwd4+p67i8nOAQYH3SN2LzQ5KRoIz
PBFU+sfyLwwk41wf7wULstdcn6GA9ZO/j0DVF7QEE5USbAGANEmpXifYkZTltsBC9lE6/fA0IK6j
a4wl0Dy14IxN7GmfY3LnwUv1xxkpjCULclYEN1dZwMQvsXJTqN/TWjUboAArpo39YcX1Ptfg15pF
IW2nzQdgIS75qSlSWTXN0FhZcH4wXDOW5eEBTSo6lwHYBsXE3aiPZtXO18Q9zTqlmlj57ipeGYtD
WZ9F3od3ksmAi+1aZ70meb3iGzVBpsb5yT40K8hKtOdw7JvFI1a5PIXUrtY2bsScFtIEQDLFstUZ
6yPOSNMbxL+1hYjPvAoKQylCX5CiXSjkIC44KiSr/I0s/j66+jzCnSpDZH+cJ2KoVSpbW4gdkquL
g8KubmSM4bVmiLHOdOy6likpli9eura1zAeX3luhvoGA0EOLAZcBniV6OWOPw5lA9plw2qq2XsF9
arjewDs+/mGDwdx07pQ2Xu0R0pcPVeFe5BYS/mxEP4wm4ENwOxVsVfLS01qN9TwrCXUBm14a7E5D
SadzgXy9m6KSgL2GFuEiXPUbGD2faoJ2mcEOfM0J4cTOkz1UpQo3mmnI1nydAjuzJ1eXBBhN9iC4
RBfnYDLuCsk/wJvTcY76CUmSn88AnJw/eP7uZYXyXMGHHekZ/pn4rKejNt0xSOedR6hKV2zhc3z0
tNeSzXknHuuC7xRQfTEVTtw/aTCzeRAmNtLn7hhcbOc91QLOLY21vTEPhWK9MjO1qSQSS1U2s3so
EC3dS98swHN1RH8zZ1m0lQjMPJ6AdwDkMCINZ8ipaLxdLLPMGOT23e8+0CsMrwnKVzS9flxPBl9s
u9s1O3dmJX979r1GaaskZWaHCJKgaXxIVrALRcrG6ycMumlMuX2R4MsSxiYGn76T7XX3RHRlXYhs
fIqQu1MYx0QUFmlSmg==
`protect end_protected
