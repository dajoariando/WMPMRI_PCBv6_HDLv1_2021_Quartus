-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
hZkXDmZwYh7Ny8Un4f/Mje7gOyts/hJRIMVKJhDbNA/TVSm+nuqj7lxONnEKp9KEmXHvp3tj/npM
ln5Ubv+AkfNZLQ+jMr+VxqGWDZ6gC8Va5Etzy2ByiLEgEH0p40N9agrHb97oD8wgMqXdKbLVpytT
SPuRjxAy2ZCYp2NKQ3m3iuNaqOzpZzb/tppBqkLYKR2ozL54KgJNACcS1bpyzP5bDX4BGz9GznuR
i1JLIn1HkoEVTjNI1jTUX7yywBfMPi3btEU+SKnFvmFIBREqh18r5k2CFOW3mcgKXb82TKj8qas3
2TS8fVMuchQ0tECETwaHMDm0lTW4CgkhyLJdhw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 45120)
`protect data_block
CXPk+yhoU9B326YdIV3sMSG3LFO1WhxJBdpOvEb0mN06E0hKXkPOxe1s1VKbIKceWnSUUvpEuxrv
C1AsBhb9Nq8bk9nS7OFUZ0jSIBP51v3eT2jzJvHrfh0fDTWAJIbyB2UVkrkV52r/TyuP4zoRpXK9
5fQyiqYklFBXz7AAcoDHsfFPdWkDNytsBl+umKGfKnzwiZE2caI8fZRan3ExTQVQMbNOA7lpm7Rz
+FwHgyZQtCMMNgIoclOsmyvTkxa1XkMBW7dKBpj9EKbzJTPSiEwoXkw84ufKI9lyMMCEIN1ljCRM
hiKQlQYJksOQbNiCz/Cfo5Q/j3yQWqrlyZb2WPTEqJ3ZC2J/W4LmdjGg7tzQpr8XuPnrs6VsFSJN
zC+u8UT/UdH0HNKWM/YvdBkLHF1o5g5cTQ+4TDamz9U4fYtNdD57h9zGLKey6gxtf5UzK1vNlAuv
9uakdy1PVmEI6nRf3uRvec+lZbEt7EpVbGC5NFNwoaPVJAUTnuroTeU9MhEmS/0e7U7Xu6OsQp2w
9Ye+3eR/jRsqznbemk8Mlv8UKJxjkjcJo6vVAdo9/3znLsDVZuI2x5mV4Z0T+k7vrFLn6stbVEU+
tg17xUEYAFYho9BrYZ5cy66KL/qAL23hIYowalEK8e7u1crcoz3GnTqkEIZB7tEAlCv9Hw68yz2v
1g2M8YGiW+KB7XFqWe6vnrMMXlCzA6xsMC51nnlRDcZvo3qBWAZdsTJ+8sWF2uV6s1jLpq2C161L
kZgx+7aU19exbyWMiIvZYjRiE9jQ/zEH78xx1/h8X0w3cUBb2DnHMWwlawuR7CtPZOTIXmtxhbMQ
kvsCjT8lRYBCCsCEKe6RLi3kQqbcZatYwKqBpLrXVg5QhlK07YVWLIEAoM2Ak303p0bBS1UfjDDS
oRkx4eXe+MMqJ6M858JRD2vTcTOpspTIu6S68ihauyIBFJ9roBMbGVjFFn5ceYXm47xf+NokKKDT
VOf150XiXMUMZfcP6xRnPBNFItVIaR+qVSPGW9d5OIg3es+wBkIKSsWYtwvJKug0pyWSEt06asW2
7aD+xxaQwlIU658fu4RV6WAd5TpEGIKyTmcmpayNE4lWyeWahC6YN8dnF1X4x0VJAheETCbY7wtL
pBIXVm1WX0hzgSW1E9U9BWOptonTmWCDnSPe/p3b9rZVrGwgQlvehxZjShZ17kINMzEqOZAhcS+1
xz8O9YAQ3i8S3JC4koPgHHus3EVB9OWkF+7afzgnlFDwDs+YWXMjEcVT1rWDUEUe2TDd/Lf7Vxgh
s2R183SejUU/JEF+fxwBLzd27JX1lmscT82gdLlVBFx6HKV8kwJ4CiQ74hVBoZOozL4fVDHxihSz
y6qQT9F9/dOnaMxOMQBcmGJS2yswgLz2fTuN9u0yvq08pkHpOtbrCJq3+FrTaBUfzlu/TU0CiCh0
XTbpkKYE68kSmUY8b2W7AHoWuDHTK047yTlv3IVkrah4At7JOJMMyVdiiNWh1jB4zXq7IOLmReAU
GfftJXGX0KLLQRAa8A6UIPMtZZyEQoU0JgVCduLRVDNhMj5xF8cA5vMh2fn8IXSvS7l5iO6412o5
MBp22UDW6mjUx4xs+Bszh1CSI5ADWMuwOba300DqXww3bBHvR1405WCk1W4J1N4WXyOd+r3PwFBB
Z12F5dJ2eaXHDEl7dx14Mn2YbWxmsO++ds0cyMghLsK3e4+MuNGJGmkEP7ISlmU4FsSduvi3Dfqw
3Ig9RgDXw12YYoDa17CfUm0+C1azfE6dkVanaSnvP318oHdqEVfiALMAWGHE1s/+IKWfMzccF0uN
iuyB6EPfB8QgkLLlDmqJzAfa0VuAs7szk4zDn9YYKhRtAoi8tdJXouV7K3PdqEtLlJxn59Vvsgt4
WP0PPuY8yUoVc79no/kAVtT6v3awvAAh2dB44T6Fix1bPPtqNp5REoUnxUdpvMVU6vAJ/w6TqLgL
K3UzXIwLLFrWiKsP1HJ81IlWxJxY8i98jcYiNqU2GMMw82GjhfNS/gdXAhNiIPqQiIMj48i7l/oJ
9u62+rDamy8uWMVtQXBI67N76E2SBXqW1/0u6R5LiezXYfmuZX5TtEfwhwo0k9IcSSOLaLMwyS1z
aFrycdLZPo0CnbdW34R8JpSAUyWGeK1i3cbkzhq2DB/OayYcD830Puzz44c8e2IaZ5b65aDfdX6F
dUnq0em3i7jfkPRXGR59OlI/K9hyqLKkoBFaciemdtv5g4W22EhrpfufM1f0A4kdXQdKJyOS8mLV
ZcYW3kGlrF1VbOCPEFqoEWXGZrr2dNrlp0Pzei7BYzY82qndYHjV0Zp7wG9Z3oay3YIHpl/l8bUH
dUcFxW4VpIDJi6afJ3LQ3jIyiiACrijaxnkVZYQ3Y3BZCXxi3cnldstFI+x0Wmkqe/l9G4gLi4AW
YKiBBrXDOvjFvXKZSU9ofljop/9lPNUbDPttLdYMvYjRLxml0GxAAsqRa0ptc0nfPqfQOIRMTyu5
XeQBJw33+VAT3B9WvYoWMOtGeOcFeUvme6MyydAn1UDyTvlaSaV8Hc4L09hWijxEBzbHMTucWubv
vltX8GKqOXovNRYWpKhlzIpJWhKnfNawqVYCe2TWtGcRbagaDgepTVGF5rggeZQv5RcUnJtqUmQm
JQG+nrpYuxrcTjojmYleBwMbZi9cUqX+sDC8buazPFuXPvDIx7GUGDRlSrssY/MniuANZzX1P/rX
oTzjqcmfUm3unVafnnK145oaXnJ2+hIQfiqYgyh7YcBvj2QuZxjLNzL/tQLGmXZ9tKg0ElrVi7Ev
0OOHjwV1ZtTIInrxPFxNwbRbv0h1DIMzmjuzH8pZXJA7ndMviEMwv8/faB0FIe+dYHijxgj1awex
jbkVS0xg5UcEZZuxnp6lcZ3rXvoS2jm5QkdHD3NPbj2u4yAhRf3iqxZF7++HK+GfPP7e7zyl8w7Z
9tw70m3/X+Ytgl0m2LypQIi/Jy769SDTrDmdSjUqvTpmqpWQ6OKO2+E9YlKs5sXglVzf7L50uWER
jrE7XJ5ENDY0juRHgHwjEV7LabvAu9+IVeJ/mLPcqwqgYJgjxWY84BIJxXaC9NT5KRktZePpPVbt
xnWsWCu1ohsrMgtFlwsD/kj4L+Wo/4B+auZLaq11EghuzuP5eG2gk/vNurg9LW8mJToYgzs569AE
jUWXAtyC1mwFEoYNGGIyIs4XrDJq8AtPaKxbq0L8CGePMTrbNIVdz705FmHjiN4EAgY+JKdm/RAI
JVTHRScWw4ijK38xr7vAxTXrv8MUnxgBmo2v/K4qImf+c+O/J9Q3YhlXfce8klomdliuHiQBSc2u
W1vj4rDoYti1VBE3Dfp/qopzczivKrTGy6Ijt94TIufxvFHIrYl8xLJ+OT95Ua8RNlsAf9wjiqDP
3LSLAfmKQ+cYpaHDM0/J/iPkg4G3VbNVazOF+IqCAp+v2jS9vv/VAAHnqwTrE+04tgqu0YLC7upE
PUfDjdYryhHI0vFO0kdklUPLPherQvO9MNT7sd3Vc+B+OgFYwXkRYOIs9BHVGeAU5t8ScG+88xIu
EZAV6oTLVxiKlirbtEornBcV90K50Cg3ue7g4XpUMLSFQXl0JjXpGlaoUyqclCBFR8oqDyhXTkaW
swWlAahvo9As3LHhvB6Lk+Aazsic4uvunADR4m6equNKXqJaGY9JI8QEIdCV6ntQcpqnsxh3iApB
b5T6XeIJYmYaZP+/cJuabMPyA7eJREue4b6Ob+EqoJsOBQFCw2qAzrGWU24iNX47KSjZJQ/hp/0W
iGyTfitGFuupTKS8BNtWEaEpJmVhhV4wnS1cyyGjmXwTgV1+vmb2FB2O7zJdT4HsfKfqHyymNSh0
V0BuJrm7ZBdTknZgacp/9lW9Okumuc6Jxl1zJJqvXreAgkjgzG2zt1+Rtoo/99TUqtH7A7jXTqwC
ymVFRBoGhEoRY8cQd3sN6S2KpQHn4h6Q1InjStWeFU6WT+gB40TIlIKYmokh5VRtnvAI6Omyo5NK
SG6j9bvTBJGJpSY8kBGnGR/tbn0cc96FUzDRcbafKzSUWXJjjBt5m8EohGpFuQq4TjHCsGvvtLWm
KOlTDjZjx8g9mg2I9F0UFXjKoautQ1HSOtw2sJ2922eWOuxawCz7EkQhL6gky2KS35FI9SNCPcBx
j0jNj7cyXmZEEEwdxQc7jOHUuC7i/Em4i7cTsAdvkRDMAu+1A89TAwqz+yG17O2qDBDm9meW+0ww
OpnJwCzyPye9wYlKspIe3LxdPk4gkAsN28YniZs/HWUpkdp8Qg07NnqzpaTJz2vmK27OURN4jyEJ
eTPS9Rf9hVvW6xw7yQbEG6jaWysWJi0Pwmv/zNxcirWIXzswmTuFBQLyXlVqpT7z3cifoL1dusPr
+bbJ2Uq4xSGoC5eGX7DrQm2DQq2Ec2S1ii09U4JqOS2pDT/BPo7adafPkWrOmI6LZ+V3ZBji1CAe
jUdyB4JDYhnsm0w7LXOf2TD40cUp/FTzN4OkuQ/J7CXiycBZlBuphGjc/HyuwdQuVI4dSSnRnjM+
X0MAMKp9QOEKZ7d0jgCU3hOf2gXcSy3rVpbmC7D3GlRjkfFoQ0v3dYIe+hhdktIScDmsBISlwI6V
JmCcNCYZ0PCbaw4RLvAFhVw8rM3OhwAzh88IqNfF1n/0dcofnMrautmO+UbbZEW8DfruYqZBg4xb
9dwQggCIqKrHAN2kFeEGbp1Mqwonq7GZJsq/ft3hWPKNH/aUl4GnCYO3uDJjvzzvxA5dHP+0GUm5
B2jbbVzw7kkyJ4GBG/+1jeZxEnLmNJaGdhWl65Sf6mdaf6Ifn31HgtinaWnR2YX+C9/M95x21TAq
1eawpPQHjnZZ7fR7WtKqJVhIpLsdMOl18lMkh0H9Fx9A+xRNfnQSHDUPU5QJomjeJRAc8SImuj/5
iOIMGScYzty23l1KhCxRBA4TkodeAp4GDZgPeKPqlGCmXTiWdqen9tIbE7oeYzmu1sfaY7Cu0pO7
Qm/cDsqZCW6GB3PrbSzxvqtKFGnDUKmwqEC4sSbx1120+xPawJ12c7TvxOK7FAFT23PRXefqzRSs
Wxsxfa2feGfurQEk2ZLvfIB+wokf2cIibdWmFBMe+pzomFQ5VxSJhMjUrf5LKGN75PCJZI8KZ019
xA9QfI7VTm2oucUDyaUGIgQcpzvs+BDzer8pXsysryFSs4IW8y0YMzx8FgngNtdyN4T79tml+Xni
64WjViNIZfNhyz/X7Rg+hzVFIpdCVJyeKT8O1CYSe1Lzp9q5oh5iT2Q7p1cgKUc3XQk8famg74B4
UrAzTLjYDFiabuGhqcBOY/Zj1WCsQ2lexLgL0wFUq9udRw5GUsty+qkp0YSps203HeY+R7sHQW9t
t+6Xo8kcrUht5qor2clNuq8NMDJp7/aB8FjJcQVVDNHcSjYKIejVY4+wALhO7peav0FKf54YnkpG
CcWDyr4uS6v9cfWd7aO5UNHMPZnAhou+doTLo0bn3Y7smf5Elc4DsaQQSowiZBTMupCQ34giojrl
6kF3mUyMqGjhYqJzhWUk5KJbZS+uaquL0sYPCFn4SdM/3A+yqr9/JOs1OfYczFUtEkj5Ov/VVNLG
DoFbMLrZPTMzFJhUL57+H/x9cORZcK9M3yBQTyfipg1q30VMZuUE0wfbH3f1UzvBPa9oo804xwxl
uxMuOsADOTaoZVbau3n6TCPPOVWdaNm2WF63NrWlahd7I4pBIUzZn1aL58Hw8JeT/hF5Pmdh5wZw
7CI/Z+i7mMVx481XLMM1nnA0G78d00lwnEc8Ay38y5J0yKk5g0TaoFhCsRtUS3cjoRXzPeEBfhf4
VJjzIAm2EW0kVVaw6Cj4SyhYp0d7xUHZLKgVUSnbdoAr/DLS9Louh1Kg/IredRrJsGWp594Klldz
T2ZvWmRjXAwqxdXvPpMM8l46D2DbiT9qCEcEByj6PRElm0tIgJmgfzPhlR6HO5NkRqWb2cPzC+6Q
1Xlbf7zVk78CTiKDIh2NCozLVH3E83BAM6r9BWLhMnI+UtTsotLiPcJDQCsmuP/B9lK7SnXue9n1
cSFUeM8u6zzIA7Kj6O3rctcWzZEniLW792OKDrb9fdJ9NrE61s/AA4vnABQxDv9NfD/mEdtq8JW+
wUVNirOT/ddyeDlhKckijrhL8LG9uM/yyU847ZiWChcmGNkicbOIeD7HBcuj8WWD7kYf8/7pNsbt
GLHn5xL+iX/56MQRTyls881pwDool2yXGbBD6de8tE/M12ZE2vfStQ1GSRVEc3REcbDlSs60m83h
gtnBusmPwL9+D/Qy1qDoOgWNVRo9gZuK0qPanMy/EblnCVegauBbOve5thnuug17z7DFO7wV7Jm3
1itPfloBYTRu1otT3C4gU2ZHBu8m7PLagOXIGisAgZfnAJBsaOqt5NeHcqvgKGN0/ywSlXAIiDK2
+RC49ID9SNS8yWx8mYxMZgAxalgNkqvHniQOj/zIKmmXx4IbO6mrgQLe/0wrQ8DmY29KdxP/W5gX
PiuSmpJAEBzeOL1d0xCiBMylntZXeF8/aJw4BCOtJaYmM/zf6v6wmLXLLwq0oaxYiK0nOlEJeLLz
opEvigoniOaf9RO0jk+Id141y3d+Si8kJMY/UHU7YKD5uzyt9SM7V/rHh/ej1yn3NJ/pHY4G3W6W
7O0871nmKjAhUOJTxtOOGXhQTBhtb6+q04YP4TvZte2W1X+2+upfUYRm98yd3/uEXe/N5qLb5uid
wVys5Rqq6e7nwD7J7kkEJEDqHdhVmrZ7dwWp5mZ6iSCFSzYbR55w6RqTnIR+dqgM7PPvpJFXLHzP
50S7hyrj58ZUKob5AYTPqz8/8K1mq2Zyaq8v4qmD2nfITahgiqurrO7RZbXCjSqIako+7Bvuvc2j
vyp0VN6/hA4U/Hy4pz3AIKsFwcSTpPKMLFI+hIaUDcxBk/8YyaySn1yhp30f9PkWVMXS2bSLgenp
0ai3gSQ2qeGv2+crb2FGLJV8B5U/Ld6cKXNL8eYSGL7Hnc9VMyQs0F1vp8Ibj8YRJQT6YXySud0e
M0YJGHqBqFoVT/11JXh4WQ3oFEZz2VSwdBn6T4PRNKyckY+5BZGj0DsFbW8U63mz+v2QIiocdSxY
tkv8ZhpjaYR/A54lRa1XiW1NoBtR/ttyYRucuSYUAAuGA+QNkxnl90NiLVqLT24OE/AHo0yeCLpn
seIQi/c6s8SW34z1Nc4X5yp/6W9wCMmSMb1vxUvfO3gtqHJuzd64Vf6bB7oBV2Fc8G+ZWrGz6RIy
gXdBypelrQfcF7dtyOOLPLNzaN39h2eK9t+sMKy4ptrmY5A2jgKPcBtYMPdayP5s5UEime0DgYrc
QP0wCGntbf18lr45LcD5VwYQb2mqeX9yxj6F7QiOoj4huWtc9j458BFzLX55VyrxabFFXhbVRtCp
z1iDooZV8fgD/08ZAfNc1D+lf2OEG8ismH9d9X18GCraoSEExqY3gq12Fq6sd3ud47+m8UuZyNjh
bVqcEGLZtSYyxiMg9bq5tXEEqjgPHiQ4tZK3zDtyK2nLQ5n0d5P2sRGjZ3JkfPjzLLmXi0u2mVcv
5YiGwaIxwOULaB+Yx3Q7IZ+jnWOj0GNxKxxymqpPa5N3DKEkTqZchj2Uzti83YOliRW/WMKBLjta
YIaT9X1tmp7C+Rs3BXwzxrMIcoKwC5C1iAsI9ilm27Po9Zt27wYOkehBHcgjLWk2u/qnq7gUY3I5
WMSJixusiMNBsheWpUQrPUUOnv+qexqCEHWR35K3Y2zI7DODooztw0Cbt2ZYPoHjeHKyJ1sVbyl1
v3KM+fc0MosSGoylmyXb9dE8iekKrgbzju8FUh0rmjFnldzkwATiE7B3EOVj4cBoi5vFDB//Kwsa
aeesV8kwfFBlmpHSeDMCyZsqKTrCA49P+mODSkSY6yRd/H1xyAmf5wT2UQPsk9TMVMCMHFdfLFqv
EFJw8cnWlaHP7kJ5SR95THokWfujoiRDTcryNUx+kdWyA4RPShVpH9eF0Rz53EEPFjAOt75/r1Ue
cr082MgUYWrLxqId1aB1CpZ1KKCYSbDdd2e+3t0RUzuUbdAHeRUF6FSM03FkZEo4ejoQMt4VTr+a
slgza6XJeIDJLKPbCMYvo8U4hSvaE0J0E5DOYAaDQc5/H+kkFyx+uNs8uEpD6gh2RgjO/83GjcQe
PC46Q/BdNOL8GE9yfLsjykRdwzVJIht0mnqsNEsD195T775DAVVhbUy9rh9lctptBwiOozzf3xgG
NzDnK/78QHtb6H6oHZ8NybicsRPkAdmnS8Cm0OGhnA0T0dY8nGqmsW76QBOqlWi+jWjBLZeOLvjM
R1sgJTwC0iWIF3kOpjNjTRffhSA484a/lyarpAkIgYDlw7kwBJydDl/BLa/VJaeN86vdyA3OFMH2
9bU9Z81/Jad/a9pgyOpGP+lvAeX65lBdTLqoppb9gozxXMetx2vUiip+YHZber6bF0TYKaGviKyJ
WEWsQUATsJPq2rZh/M2BLJg3L/PPwnUkFDc/JkvIzimddb8j2nykkBSM8zwwF66w3nay+IBKwUbX
GhqTG3YfemC7Rv8/ski6nyjINK18JIEWFoY1oLHekYCvf6huvX9kON5Qq/33wpONtK46M0wzYxwK
c1nP5MP3QHv6KA1KVVNUI7WRwJ4JZaOBv3B70OJVVSAa/i9O5U1umUMYMbuZo8rRLAqIHS3368T0
IDuRYNRVlX/FsSbNJcdo5YO4XbTACrCFuW5tdNYYNz5etLYibWKCgznkrQSh0y6Pzvgv9C1YA5JF
Or/hzw0kTJAq3qzGdJ5yCEJRoXPSUPC5mlc/cisJi8NUqjOc1aSplODZMVexyc4Yhu+Y+4neYyRA
GIf9dhqfNQ9EUCVKQMxDnxnj6pn+eVH6As4O+Bw8s0tVH+L2a+inrWXpxvmBNfmJlOsMfu7TIZJL
OlJouG/10Ti4fCwRkJgFfoeRARaY7k3PiULU94Y0HGkjszko9psj0oKbbx3AVoC2neTiyXpDhs7e
DIwwYL+Ka0iKS4D5JU7PchJrYUry0GJgX/pkYtCOwFd9hVRShsQ+VSMB6eBZQdkKUNbY3wo2I0YY
7lhzW7cDJvdJG1DGqd2TpIRqC0GUDJejMKUHCf6L2Nm/4fWXnjNkpbb04aini3SEXOb5yyMJ7IXd
ipzWUN+bNhYj2JO0029uSG7abBsfzsD1D35/eWCqWx/kg52WjySSxVnE/AYoJ1JmLk/EmjSqN3hS
bLn8AmDAisT4MTSuijb6mNMiWrXVnk2ElN6DIp1luctetyDI//fgK7MnwHvfjmljsu+r9IGQ6bJk
R9NY6fiAZBfODdIvogb8PsoC87/eJL3CH5x1wDxIRXBOd8NaYtkQuodaWDkPGjSDs01WMx+ZFUQx
c0jiB/4IO6hcOcQbF16dOYluceNmwZq74lA4BLYhwvjdoBlTNH2WmWikgI52oWwIbnB1SBKRmcdz
8ZXw+KGLdzytZKB791Gy5znCcVBF6zPdwlKhJb2d0L4aqK1/k4hfPfXfPlMz+idtzxgrcOJnz0rC
xNvsClSNH719RnAqVzr14ojn25If7sY+5+x8oqSP312yeJGqGJhCGLu1IZ8r1+q5H4fG6cuPaIhp
B4JAV66vgIdm6xBJp1LPZWpLZuYFip0V8NDF6ZEhesYj5W7xVWnUehRtorfMgkaPZ03iyWT+4W2M
H+NWjXmW+2oQXZmBkJe/BXt5LTvTp4C8FKasKrDXiHGcI/qUKXsMqJ/MxMWtIPsh000/AT7uFCUO
H250jMO1OQxSJOBmEZh7I7E7WZ8EaA3vTj2BRXJ67tpvX95RtfCzXWxabURt75BSO1wBrHcqzTaK
buxcXlwqYa1L8BfIZv65Sl5yhcEA7xdOFyRfrRgVi3+3BZOcOqMl2IQOiqRXSiQrGT0yozVGbfOD
ZvgyhRFkalYqBx/pk/MGBy+Zm2qvApwEmAJMHA5UJBQ9kPtlzugmIUUQ3ZNfvps7ACqPsvG7GeW7
SEpW+JTb1WHxlf4y+ri2TczLcHjP/sT1YrLysPXBa3SANdg+TgF/o0dTyotWrBd65rK/aqR9KUYe
j/g8wkGf5DtX36cg6VwZNWEt8sBxtzSjjEatYo0H0fWgmT8nz2lnz9y+zf8dpwk+Eu0hOL5CBJxo
9WnrwJVnZBqx2NAAH2CR7dY+2gD1+mt6bFxH3Xh+brYnIo7nonkirhov7b6aoy6gcK9YyfbukmyM
F0suK0gHdwyEqeMfJE8pzyr4yhAEP9tKyUAVpM8SSCo+jNfHLhFQYi5lriXTA7EVkuYdwbRiCpKZ
uEYm3KOgP6DvrHcMEWIGrVXT+ZagG5qQheh6S7etU/wDs9iNgIyyt6dlnb/rn/qDp8qZXFNRuW4C
Is93MFPYWQV7BU/9LJDpNtPDpc9NfPTzOWAjv3pQc8TD11EH3JB+BkQFv9X/Jo2qxCBcFw+SZvQH
bqxNnfhhhlPl1wf4qlgjK5RPF3NCymUtgDTXn+Luytwkf7VCeMZr7tMewiwl5jgMwj6vG7OwPsGq
u29IYPWNr0CAlsfo3PDtmAlSK/X2Ie0+77Gc4OoQVCbf3gUlc5Ifya1AHqsIKzCHvJEIJy3g9gO3
1cjStxMA8hMRZCamyG542TvrReut7Z9O5968telLwWd2aEx+JImhHE97yMvRDkvD2saIWs76wA1D
xniW+ekKJUxpQvDt9XgIKmpWxThvhu6fC6+dUIdqUz3qr1fSD83G6NNzaJ5U12h9waKneEescd+n
7aSEynRipA4zU0fcX9REm/u94BzL/WALjkCoUhTQWqy0juiug12cjgsIHWy3qBzKOAzEx8eDXwC8
Q5v53gvDIEENMzIyTHI7+Edc9Ry9IyCTqK013FcOfk6+a7U3d3J230LxHYnnXhw45ZvylfENiDB+
3AqzDFLABSkp4k2o0gVTY9/MuqjHV3+PWBpQ7HqwGrqx/sGbtDUvuRP79AeL7h38NmJ2Uwx24mCS
RJxD7Xld0fUXIJ589SwGfMHuDCdfPQpXoBeqw+l7STMUr8Rr6CcZOuJ3uCvqWN4OlRD1ODtGTSxg
OBOsS+J6QelGrU7jXkDLP11qyROZ2qFsMu4UwHxxR033Dtnss4hYhA0T4EE0UO8jC++SPHFlWkFt
KE6Jcbrnhor0E+qlmYvDksuTTBpB087W2jBA/Sndinvb/09qB1xne+xMXU/Fk4AJM2vQicJqBWrT
NTSEsSUlNSQCOIj2rjr/ja+1u8Ejgnbc9ewG2pG+sJy+/C4PEf9QincC+REaKzPxepmNQitQKvNz
t9rNB1i9bnxyINVrVjhQ4RTWcWGZ88ZmTnv+oMkRFBb9M6r0jsk1erKjtdqoLs9i22+gclXodsFZ
Qbf+uvLpgKySABnFBrFNHjY5Abb/0kEBT73MAYqGL8p1jpBinHhUvH3WYv49oN7sFPleGd/m9W3g
RxwTtsNFJdaTT4rmm6Zs+DUmKCPPtCnJ3lVpp9xDa1JbKAChOHKKZd3OLBRVtMeS0yH36AsK4hvw
n30y9aMzgp/wPbpFpgS7NN9B4WWST8FVaM5vfmSaNYJD08GH8WTD+ZsLor08n/W7ZXTEJq5OaG4z
vOH5Cfv+ZP4eNKxtAoVIyWnHC+CvmYIG3UrnpjlKD0+90kRgqnLk7LwlSC6DMhta0T0J6uWjgRD3
JGvKnsDpswsxSGcuHhslwCFlLwrVFqkkGFIHLSea1iQNYATsibIbMGNj7zXzjduyRpvxZE5nCulE
prYuRvLOqL11J5MHBtQVG+5myqJOytYJeZ+cAdryGEtEO16QoRNG3bIOFl9k5LRgGiM+7GZ6J2Qm
aV812C1CbfqMn6zIFWLax9DHjhHdyXSCDcfCYQBiW2nzB161ENKR24Py5ynLz3A4WPl1yC7PW0EP
N6YfhokHAhWr6RKTacujm6V7GwCYxsnOwSPW83YECjnX9KD8Qhy6szVdn6h6avEbCS4DhPokhYHz
8IsglPf+CdfdhVDlLMHNi3zVkCdKc4xxCfUC+tD11laySlmyp2pctSKO3Ju59wY3Oe394/ZAam2u
C3Fag7pAWDDrdDdXJZAfigT+/yx2cYD5iQh2Jic82zRi1A5kzF0OFOkH99Td5HBrodtZt/XoR0eA
Og03d3i/wMrxzPDTGvZSdvPME6IjdmyNrcyHVF1q0RrfOA/2Usmxfc61YxVx91nB6jcgAUGJGSOr
q14h3XZbvPOFSBEpN1xDuyfD7S8Tgf123qZCIWQc3yYpFaaGv067pbiriiJzucKliiiF9ODQblwK
7RkYQZWc42zymY/Yzn2EJnrc4yofMNTHPNI3KiGqixZQM0nMweDNl4M7ShLc6VCjoLibAX9vuUsO
6519vNIBygt7fJmGT1z+TOV4dN3WgwZ5DNR0m15bXjaoMy3JJbu9+CLI65SkgCMKL0oLSpCUS/KB
KUvCy9u4XtbiZq5zhjV/orHrq4n1YXmBifilZVopGP6xpi+8GssstvYoOTFQSJh0J92QZstGp4Ob
3034tap2OjnFidb9a4+txfz9vklq5WmRsM3MvLXQ0TvuD6uIYROJ85UBMIbbJJ7IP6T0Ddqiyf6u
6ubSD7W5rqUC4EwR22s6dIgYJbqossTx2Py16gn1QgW0YRyBQj5XZld2pixAmNpesGRSVc+dmGPj
c8ly3dU8n5xVZSwD4okaiyPolU601W0Sa4SFMHatNf4JhoPD0j9IJhBBDe+ZNeCXYh4Up1ZtzH5b
tHaXJ4suhCZemkB/oZzYcnehA3JzoMDDiq/g4XIGFLwuPhHcqmc/4Xe7MhbfA14oXLpbcEqI0OVB
bere8yr73VHODOd1uziV7ykoN0oRvqwfUbUwCHsBcGilHie8wkWmKJo7ZCkLTKwQ21TAwdFvuaio
9vcJr/+g69F35ZS6COpWzd9Nvs6zBEAAAhknafMKixAJzJsAtY01AlcvKtPZH2mqN/LSs/CEHDZ3
8qiifYIGjDE/6NFNQvz69dFHRbA5/qV6y9g+vsaono2Tzyi7E6o8x2L00daydYOKoVp/XPv5zCpN
rDH4/sT6QtL6hMVhe/lyEDIyoEBoo+Avwq7Bq+mNc0SstMnb2kiEa7XaB0Oh+u1QzluPCUyEWh7g
C9kRBSIsse5AwsdkTNyzwV128YbJaeKAG06ou3YPxr0APE026SpCPWVp5n8T8iWK7hkSePm8Vvo2
5EtAfASO1ry5eVM8lDWHxjy7/OPSdxemyhHVOJO/fX5OdzLqLP76F+CDqO9HMZTFy9HFJhgetAbW
hcDBNsTdOMhQzHCF+h5PUanEdICMsroOPP+z/CUvTIx2rZXIUA41vsXWWLqHy2qVmLd8MoCzaYwY
mx/bmOQqcLaJDBgtoQnNKtIQDJnqMGW4Zr3eYaFpptyMY6PaqnirkCKI51yOekeNe+jd0Mbr5DwX
O5osDISo65SK+IjdBdxO39avXDMUx31Mzbzs5WyUV96PPrrblD/OqQRyic9CZm2PnjkdYQFgBgUh
vrurmfmnhkDDFd9q4hNL1RP2IBzLuBWK7NxfuvbDKIwn+DXDDxmpAt0h6V4CNTZlwl/ZiYpYXJ1O
zmCm6bm/Ars4A6NylPUb10FqyDtpJFW/sprz9Bpm2MkPwDz+0JkQBGa5lC07fX3+U0jggiEj7bKG
+frSfFcj0/KRhLdJwwHnkl64D4pRUBCGy6jlN+MWgdGaOWQAHB3KHuUa6g7kqBaZLBmHYYSrcDDw
0adMy10Jj635m8xsbP6TJoctmtdBMjiihpYRPvNsuf82JNy8vUiUcG+R+m/52EFM6ep/KAZI1zb9
+jLZANsZ9HCPCJVCrm95QpLVrH7aIsTnhJyYHVXpU6hZ0NEV2yhhGXmPF8Z9SHn6rkv31AQwiJJ+
mXQX9uCP0L5D7fJVHOr3iekwJamdq8rwiHpSyZqXRVBOWVpiWwS36k2er1+UTmA231QV3mwfk5nd
XpFPFH9S1eUTSe1jMVqSCigbqlv7gRsSXzE762pUNZqufl+Elh6V7zRZVMGEwCvGaJ0gazkmAZO/
/xLj/MuzRsMMF9vbMp+UExn1X94NnMLLh9G5bMEQmblP6ZFdNbMQq6SM9pIbfho2S7FymmaurrXn
dYIDaSjY7sDL2CnifEUCEamc8VHKx/QtN0KDQ/SbHBge4F67Ult2s61HuqVbXuJkmkAMRdTMGpTd
/H9xWsLx7Tuw4WCymOBEWFRBs6oVtAMjrntDx4JqcX2kRsgbgXVJ/LY3ADr1tOJ7t42/vX+hj+mN
ARrUmSi12HD2Ea94zLxeX4rxu1d0Zg6dHI8FgGgwM7pUxOiRs+utgDLibTRMG9+YBMDNRrGblzSA
3Lo6zCSOeTZzqJ8fcgc62nSShkU0jISFW+qiduJCEB//a015Y4ZCo4X4LYywfBhCIOP87eSOWbz3
HrMrD02xqzzxZjzXoR8fZra0GLBZXNT0jlJ8Mlu1J8ruTo9uUv+2y6/C0+P9UVW+vqS3Dh/xpCOn
rMZmx4fWJgiFWkxJyeRXJWeL41PqQp7DTUzlzMXwws8CgLkkjFX8jjHbke8wmVA+z4d6Zbq9Jao+
1z5u6onrKeOcRzTO15zOx/ezUBz1lR3zw+lGUtPAgXiBT9nxGtW0qI0xxuEvfAzggij10izKwLLL
SxqNPaAh15JuuCQ15Q+LWBdMM/fCKd6X3b2xE3YPmCo2FUZNij3aXQ4p5yaFL3JtaJm13U2TIN+E
zcVkuxNw7GJegD7e9dT9wb8b6kNsAHjknxmI+4dOWRI/e9UJi5YQ9vH8fWCtqLGxkBtbiN3eg6+K
GCSbXOdU5j3xIeW76kEH0zJnD06+4UQ6KcYfNQZXUGV7F6xHiwSaSQntL4fOqFL+pcWJqWflvIn/
nbAV2LbfziH00oTsbMj1Lyg/M5NSGLtvjZZCR27CvXlEJPKBDAbTEJbz178m4hIiFBCACmjw0dUh
T8+yLmT+RjcmpHl4YLlynl5Dz0COvRY413zXAOC7BCRUyz/OubkMSpnWLZlsqCnUdPj1hq0AfibY
+3ZsROrABjrWH+1rv7n5w+EMwzLEY97iCDW39qJmOIL2RpVkLXKjbl2mcnQPNLxoL9iTny/RVgJl
4lqw1GQKVs2Vh/NSvNnMwSHzTlqA4eOU0eP62k/cxuhXVCvryO6PDNFHqoJ4sEabsMS+9TbvaG7j
g1DVCzJAnQjos76TrCdFOTKfNPtHeopSOeIZYvQ2U4ddDlT5Ew16O9GXSkb8zvhzvADqzx2U7X5E
i/MQdsRXtNTBZejA9pN9pmbQU/fFMjjkK3+P5U3BxhQv7u9KXuPLBtzyn6fz4bOAzPvPyM+W6hrf
9KdATEWS9GH7hrO0YPW8HaiRUKurcHMluI+z97dS5K4CtAcSd4nmADeoY961QCvxN7A9kiaFcxCM
lf3ut3muwdGmLSPsGVvCzuIg/ln+Zu/qJ7ymhJUIWOudjxU7AqVb9EgsZ3FqOQWgktC2HpgfP5Mz
MpbNnZBYudNC8W+Q5ZaYqRYeFQkrijuMql9QPJKpU4kHfgMLfksQxT68aAEBY86y0Ng5lh+o+QyX
Vk2x5WJwrxd+lbI65CJR0r2Bo0IYPKp9l8KJqDkcJXWFxYBEzB4obht8us9EWYTxosaj/mA5H/Gi
IITbBQpE2RIpqGLjQ/2qLSlcnTGwbjUCH/AVvDOpARnqeHcRHnPnV/Jmslum3uobl4crGXgmPbGE
Ftrtd/AonMBHl3ObeYgXUifLLx/9c/PRupCCu43CVpCOe7j1yrVXClcVseYQ15O0vtm3IX+c2ljG
63nTp+kk5UFXFkga05IbMvSEh8x99zv4rg1XgnEU9qaiS5l/Vk06cSZuSMw+DcpaYTbIxi32c5k0
1rfAii9GMDhlSFT7LjSZrIeMqMtEOaECdfuWrHqDnKPDKJTiOEVTd8hUsshoFbg89Y6DMCq829qH
STo2UiKBeauxwV88sgCvHJzroCht9tbd0WzQmWIs+i76sV+s41+m1CdHWhfb4vKnSN33rX+gwD1o
9IBwq8skRmt497eagu2yFvmT/EwKadx9n122X2Wne3/5dWqE4C6EoRdK2LeNZRTn4W2gHPzA+6dS
KejaOvQYprG5q4Mm6Ces+tlmmxO8c5l+Fr5SCmGXnqZsJG1g02elGdajXCdxYi4WcllJi/DviwoD
0IXJgTcyfbuMAmmkkw4Hh5Df7sGhxLOgvjII9PDC0ZHBgJG6FQKeD8dP8NOjN+HkH+9auTxNigAd
4AuNxVir//uMUSe/bCs08hcNoHPT8LZzfjpjgcoq8TSoW76W7BUaHhzvQae1JhZ31aiw/zk7JIE/
GGAenpEstUD9Xd+KAqE7/roJinae50Hgpzzh2n9mWUMNClr2UOr9r2cOxVMNdzLVqqgqZKjgpinA
4UAPnBkSQAPNbmXBQq5QkwW7j8g7HUbedUqGoPmKjNfY0D8FzN5iWrMBdJwch4VZWB2Rz1LW0UzF
vsC7QdsL2YAiG++umTStkMgDxKiLIZEAsxSsuqKRil/GpOEDgLMPy/89oos6jft5kLO7EavRp/Io
TAe+QEVRA94hJybWgXuRbhHqijmMvKG3m47JBHuGb9Xgox+cJU9ANvm85lMNkXFW3rX5uBzr7z5v
6I8UvTVhNVooCBpSZ6HAxPSWII+c0KE4RXGT+fULKGXk2A8ibjEqbh5ObjAXDjM/npEKY+Nn/tRz
jxrR8tBTUaXKIPk4k/+KkkhVEvlxRRmhU8l56c9Lc8PHs+tmDLIHbNSPDxKNt1mmAfqHw6NHuSIF
ILCMCIvJI3Oq5EAwGI2smb5bSrP9kuQrDgJOfOus7c0tVfgT5n0O9ICO7c1SEfi3EkkyK9CZP/sr
HCRkDa6oOMxjrqLnxoYtmrr5xhBuOTcKlNCl2eXyw1/bhtomzu2lF7K4Vdv65X30oupcAqE6CQU/
EeJ2nDkWWxY8kL6MF8FnkYo1GfofxYP93vuEJ09VWyJrGQO62Oqvkd4MHGN1gEuBCO4FW5ordVaV
IK56FRmnSsc5Lu9nwhQf2EqNGmOpG61RL6uHUF0euPqYn1IpYtzWL/vulBBA1cnNqfuvIOM377TV
8pZ5XQoKjYOD2uUDJCvYiB9IYWMwld0SoZh/NT4RG7svPX0z8soQhuQEgeJxPMu4hCdeWkwQKkXS
rqSaKCLkzLOOXNxtvyyxT6bk435uaJOBFUzSLBssnredNqxCRernspUAb9gQuimuGw7pOipgs0gS
purkHDJrxge/luPklgOPnpa0YOlCwdfnmbSsyHzXyxjsVSiWofxEGxcOfpmI1F1xiJSYAqDHtRH3
uhYquXCWkQXJPsV7f8hB9I7UXt8a3x/qFATDWp1u9qBAfssv5MU9YmUjE+iuD6+ETGWRAYNWp5GU
ykzaPZd3JvatEwX35oeQr2mWSRcJGfnoQYC+htA73ZomHKtuf9YDviZS0yntVLxkywThDEP8X5O1
HCxPgl5YkbD7lKmDu/13frZP+sw+UjwRapJgxhzpPqwUhizH+wq4P7zxLa5S0PehjA4kKJpgYBXC
I0o9QNLGaOTI9LfWUVUvBFJiBNeYuFce6yYS8/iBTyVsdNh9aJ9ZUE/Taop1eNdFz7bWC3qWjqof
wD8S/iXeWz9LGKsRpYE9zrkhuPK1vOfGfpAdNrfU8zwbieixwH5MW0A/NG5GOwZKTa28K3y1rHCx
ScARKbxIjVOB/BfGtjQZND5m6bO78f0kIODFATqicD1PURRgcJsMoxX4/yFLn5GTwYNyPogE/TxC
MCwmCkNfEVTxvScYzHHOF5mpifPrJOZhAb7kX8HLBpYs3E+H9a5jfp6IOXYidyZvi0RxOYYDSeEK
lAlYkW86Ts9yuy5fGbkEKm3yASSYaeYNnQAz9CnSvt2rzwQTxHbRRh3auX5UfReZtKAsbpNklzCh
zDuT4QK/8SRV0J9hunzeMEFCqowIpjIKTD5nKJuCyIhfvw5aZGlvd46Ry5Rqea956c1lBQl/TvnM
HvoMviIssw77kPB5sZtijMyF//89ajsvWmdnaiHg8Xfc6Op8cHd4Fbc8usqHL+uLbgx/gadoAmqd
fN5k9Ixo2HtsoMCgUuGTGCx/WUctMBKAXJR3ykGPEX/jySsaIG+4V8OtQ39r931x+/ByTlJlfLzi
lFsonP/O/lWJe8clx6q10L0jIcrHxktdNe3YLPIpv8M4qaRsgvntZXrij+9toUmydNk9IFyFdezj
xKRP1ii5q/nVAlaQVchkiJstHCP8SQ7z8KZWFSOy14YLUvMddhygSntqEE+8Fj8b/CKlE9MUlXgh
amTBAjfLCM5kVjmVFQDj0VNvZsUYrKOwZy130v20p92qJ3E4kSdd2eQirntL0I8qKQIYA4uDx9ql
Y1EJD4lQ3OI/aBKfkJPVQdsl+pf0eGmOPgqUSeieuoX9O+zK1GihDHYlT0IvlysjzScRfcdGmR/h
S+qown5aif/cc5Y7f3omIlRuzNQFnlZoR957y4aJNgawWKZab1L3BeKZY/S0flRbJMzXRrnkz6cY
5MVwqzEwMUQqsOBy+V3Xu4NHLsAXaJGSTWVbDLh19ajUjbxQ/Jd6ZGcgCbXEhYTAY1KPpwsNr/lG
v6dMNU69VAvAEJ4IM+LfZl4bLlQuTH0FvlkishYrwi0S5knKrTNcd16UdzorNk9lPYFGv8ua4jl/
VSgfdmLnzKKofHLFsBjskNSKWeQybqNVjXO7/UOZQBj/Z7nmIEEl2Df2NEETsuTMTboczq4ZGTAs
qtJraUNxOwsl4zJPoFao5t4wHryL2sjcACx88hemOkreWLHSEOXnEO6u7vY2G1R1dikbV+Y1r8Z8
c18txUP9FB50VC2vNlKS33d/GoyOqNQxfXQkn86RhMRmMbYUihbNQg03asVss4GR5nhuzacFQnin
kaiJ/29REKCGdhXFi4RimKieTwu5BS9plcMmatzmhhrqsq04PXSHdLj0BqoqwyN97b2sTAAbiG3L
XKjblUk7fd7Rrg8FMw4Vl29+XbJkmzGVxKnS6OKU5X/EkUyNsArhzY5a/BSbD6ObW9ObqBD2Vgvz
aIRxCTA0JrAndJTio0TfA1KaGKDrU0nYmttpyEV59N6mn/puVlUMJGw8T7G7WeeFwUW6hYH3P57A
eLtFLC1/CS/xjAkZ6OIClx1qrYECefZL+IdAL4YeJuvtb7aNSsGHS2K26xNfnq+gSB/p1OLdfQXi
sN3Wa6XHB9+9l+10tamwag2RxZzlZenYy8U9WzLQWbL1fQZXOwuocukRk8nSjG6sRNtLr8umU6/K
ET1Ikq880COqUvf1MqTF38hPeyiOwd9lPFERUTIyJ+d4FPu9QizhZ0MxXks82KMb1X2F9wQyzSNV
9m6QAheP0eHIqUbQd6ehhsFsbXM1v4VrNaZ0yuiDhEfpC2vCUmm9vdtfYM9I1cBihFAKaiAYp1iV
5B85meWuaQTpdrsxVpylfNctDVBqK20RzUPUXoLc0iEIDg6BdPFsINJz0PwfJAJ04uqvNErCnr+z
r6wLbzBETK0p68EpXQXR8UncnArz2YIx3pkbDW7230m139bUsVJRZjIJmX1uzZm3lEaGuvvI2HA+
O/XHVgqEnNepVbkQwNhuDOT8/z8M1AmLyZ9FTXSSdNrAnUGZO1y5teVIW1HnPoPnUnJfCczO7ZhU
Ix6Jef01m9O6EmEg2vvyFF4bsJbp+XXyBauJLLDv/WYWjUbse2GdcjW0AznznIZAGdaIbw8Ypn9v
ldcYmGdcFJLv5FUX5jovfqa3OunBwqDsutLPgJJP7kx1Ih2e4BRjZpCsS6sL2RIpwU/LChmxwozL
rsbJ5cOUsY9hc8muCmkatOObUh5ORI4U5CNrMyYyIcLZDiRkqV27Ol0rNsGoDMjGn2w6lbzzPqwA
RAvD/5YRm7+EGOrNO9kAUHd22GlFNruwW4eH0ifXYyBa9Jzp9r9JUorMeIIWcxPAS56qSeaLDEZb
ZRmapMWbbTOy1hm5U7rGtKweu1UThzO13jJoYHyIPxwrf2O13U/rFosWubgPlbUol2SsbGAI4Xmp
AIbxBpG4h9U2Wp7eZoJAeZmvIq5aY6kU44cKeJxWCejIIG6NDYmIwaZ6ktC72LpZd3ZqQsNQBvwG
71dyw7LF6xeUn+5WSZXFCbHWKYZ4qf4ewVwwrM8BAWR9mn0IlMKGtRkwGHmIg/VpfFZIt4h81+o4
pViQM+u3agW37JsjOc2P4RQ5RHMYBRi45O09kIu3lnbaf/epMpHS7qe2iHXhy+po8cGvVQvpUOGM
wRF9YH3lz0/OirUT0B5EV/DnCxT2rxfjLtFgrQ0yVvx2RsPi3u7ATD01V8O0w05uMA5OgbRqtSWL
aUTYJWPPXNiRSLJ1wnHIC62YotEQLKOWt9bE/K4wJ8DObgwg6jc/A2z/4rIfawNehrhnVaFD0d7Q
7o9/Yeugo7y04lbXJwRkLUwPwv/hHTmrHdSRHdCcw5DtSjOxEwfQt7TwOcyQX0Ey8FgfZYDEK79h
AqOPr8NXfCkkiQaD2ahRiOXls5DXKpMeVmDZmQdwOt7FT9glonSSlYbiRaWOj1hMXM68ZNBGxebF
GTMaDE8AI+QTjXov3c+kX0lZqh/qhd1QrUKRTZKQI4d5LEmN9m2z7NnUjEWswqsGXPAVbaTwkjiW
jF/PHQnrMtcf7Gke09+rY4+DXialWx21ebdjWbEz1rv/tMeU1cYOrTsznPlcsctmAgQKeEXzW70v
WgeXG/HE9lj05/zBCvVJbf6Ox+m3axmAudnEsCmpvqJ8Jlo/sIA0vzCWuPy2dMfgXrxcbOwuO/jZ
/FfnYQIsuPbyk+lViBljFEWSJkCZFRRJ7AgYONPaRblo9jXfu5nP/3NV5EtWvkHOPQErFpJI2xvs
Lf3saYvFZctS8VubYvXgX/cqWkPgI9mhKK23PZNHFaGIcTo0Hp1/r5JIx55ribUi3hLc9KqZca0H
5Qv2Qs/QdcXXbLFykNWTzGkInGqjDbTEfVnN9ycc2Kb+zKVcDdxXqyrpLYokI3gHmGdChwFmWf2g
b0hxki6JyvYfPuVQrzcbLHboOONTuEQ+YClEyTKLwGbRfidEwidM5dmbprw+AsMd9bzG0g08/i8z
XEj7P80AEyl71CtYIzUj92Hb9ObMmbhM6vF3SULP96e66BXFGuZ1v3KyDie2VNkJBVGbRf7GpryG
SBECpFCjRq8QCwYq7mxKvlvbknb29uv1zYnfP/tbZbzVeR+CnLtoDR5XOpPQEFw6Yhvx7lS3qZFI
VdjVtSHPDIeWdLNqR48rMDnHusQULvK/jKtFADk0CBZezNiuELJJRrvDpuIkQwDdxGr7GdJhxXmo
seLdxbUfgv96Yb4ATmWjPw1coHWAYkTEf52mrk7UwiWnyIPQ+7XfDmqiQZ3JqyereuZpQIzCqj2x
Xu517Z96e2Us8RHN+0QYH6T8k/fs6G5tPVKeIg140DkPIRTS7SBTdeO1qC18fz5Q9xATNjzLm8qc
sc1UBmMhT8hCXWKLSMZ4Ffq+9ohBo/5UMVUl72HDvSK9ybVT8SqQ+dtPgNJ2X01nFZkUzp2H5scH
gPQm7Ex9LbOC4HEZ7nWLVOaFgv8enALfI/pQOIn9P6PBJLGnhnYuXSkpc83UsCR2/DAm2Bm4o5CH
GRWlZLEt4jU0ye+Kb8i8b9UrhpPXShn7MV6B53sXovhXmty6lW1Pk/nOIEjLr36GRJSRDrfkj1QE
qcsxXSssI78htU2yoDHOi2v4mnr/ooIvv44GHHinjZx4UM1XctpbknycwjJ18mW7ZN6YGebf39Io
G4Xeq8nueT0GpkoGlkEC6wmrHl5RQjMiihNUGiBFsO5nuxUV2JU1DgV9ipISY/A+LLz/D9iYPbxX
KV52SzYB2iWwQUMcCoUF8GFRkmp99yAIMrJR/ulEpCTM4vcb9RwxZPpeF5B0GyRayz9HNOXMuRp3
1/cK0NzW1V4H5Jx/yeKO0EjCXQGHuIJ5DBdsimbVWzHmJWFplYEGgZrWmWUUAfutO5+bFBGUenti
qBmgt5oe97AapMsxbFz/ZQ6tCLT6zi5YsCWtYpwii64hhEHFcUcUnDFjWW24S9UZ1Zi3nswAPxRP
Sg4E7ubFHEoTHvOq1FNvv8oyBIaa/7B98yD/+/GJAD4amle4IUUimka/NO0BVLRx0YE3HBCyfMOK
g5PViK6lKYkfKMOWv/bKH7YvKAIYePgpKktgoy8f0uKgqqn6SGPt2WUawv1cRMG+pZj/o9KBbir5
AqI1loXGXjCYjkmuur48KiPpu3/5ZFZOts23MDpKfVHf3NNKFH1E/CsVNjzlJ8f1WSEjHqSgEhpE
haUpEK56wewDovmZ6KzyhsDUNpJ6lF88oRm9VU1FAzpXU/mB2Ar2gtpbvxKJOuMfAIrWesuFL2DG
pRoNOPomPttLqmO2w3LYY0jA42yYMREuRqLw6jY54cJi7qf0OJMrDrejI8PutFvRHPu+Y9cDsHRG
sGF/2eSD8IjNcmc+vS1NiUqj5WDypyG/aGjfX1Ve7b/P9aQFm/TRZDEZz3v6Bmm1osFu+LVauOeU
pckOjuh1bUK3kAD9xk50oPT8A0YzCHaVXK9HyJGCoxzt+i9RGyshjGafE5aWYbBbSm6iKk4VKupN
6z1n9gDkMgRKDu6gTcTHmDPgmEV11dlsd3N8ODoglOANW2e3iyt7hBhowCjadznI5tVIiRfQjBz0
YpvpffyJSV/wm7fZTqIA6EShyL2wousuv5+0dqvdcsI8EhAffpHzQNSECr910XsAp+Ow9fpADQA+
mtO70vRuuD/hOFTvS4E5vhEDhqVqQL4fACPp6dlmmkVeYJcjqKrN0nFIMl8sKkLtcqz1/oFkaqJp
5iDDUIB2sq9ohU2Jh/WQOSFBiXLaLbxYlYXkFWMVk0xzRURxFTAPEfAUGaM7veCcWj0N66s0uXBD
+RpwPozwuwC3VgySJLDwuh0VWeM4leAL2HhhSKW9GQ+nCSbsHwvZ1eMxwWjPOJJl7xra8lSxV4Rx
92xJ65aT1Ipmgm0hjPGul4Xy09YVwggH/28AWMlJz0yr/Cqs96ruY5/N1x0sZurOpQxoKebYSMuH
cq1xX17mNQDC+htxbwx7UwRjhuDT+taR7A+WC0P+GOdV/Nmh758bFy+Qm7D//v37PX3cqiAu3LnX
BHQrVwMQ7T71x9bn8oO//yT452VutmBGp8JM+GX/lErpQn/+gK8JfAlR7MMKqm2IDYmvb7WTa3rM
U9oH//n1xO0zAED6SyjhnVdeEyIg3MeGfi8ihBLsb6pETRthmT4uGmx+aosvRotqMx8NMXG+7qp/
BllKvSQ/jSU1kjHGxht1pEFpJI56MBsOXiz8n9i2CRladIWsYtkuuknEd5GFpmSxYm528iM6W7TT
DqwmUgrnSjFlxuMBbigq5YJbxKLyGIkgfLOi6J4VgCLLHuRvX88SvmHjHulaZMasfGHo29aAqZex
uVFTd6mpaOSCSowkAwqTuOJzc9r9NQwTZhvZxsRFNjQNXiCzm4wM2oPxRwRPH5FjoEER3uZeMvFL
a7fH/uFC4TIht2VZZNAyu5BAisynYZERztyE5qpraLN04VWqQv2MVP67jLq6kkd8PqBDeL1AOBxl
avhBpKQCHQYOwgUUtKOUmTtYVQW762Vi07DT7FGiLD5nqbbSUufRSjTGF3s07782Fhyd64JA/H7c
GBuJgMiXQVSqC2mqfU8X5RH5qbxpPHHMw5NmylIAIVb7leTWkgq3AV1OrRRwjh2ZOvNrenhinH6A
XSbIR9jjzb70pxaow5x9PHRM+fn5fvc6hvv2HH0bHUGgUsF/+xoZEG3ggMCVmKk1dBKrIhap2qgl
uQ8UT2wHuOxw7SVjQdJT52EiYPAtYgNWMcG5Io0ypmgmBWT9DCzZLNqIF+Elo0eMeaWkJjiH7IrK
4SjKHeH5vS4sbzRtRSkdF8JSRvnk4Etr8OXBgR7dO0wmduxAYzsWFY4sGQiXT7wp+pq4bmn+ikJm
nOU6qRTporqq011D/k9Dt7Kv89JXjVCbcF++eNhidYBVQsLUd/rUTIQghK3i4dbiGOA1dHPk1j5q
IOsgvQXykwFWZR6U5+W3ykEKY6dFHl6GGnHuXVmos74Nk8B6fvdxrSldC30+B3+fR4TVNmkzX8dB
2b1IS0FaMY4/kIp0z5jqY22rBkn2yey3QnBqrll92b65kUECDwJ219fVf+KFb/oR92mSA6Ai89dm
BOpCykjVCO3pi7VTERkgHwDblfQ8w5TSAM9fUr8H23C7p+LwdsIUKPT5Xat43QaJJGcLCpE5gDbf
02rXpWQAKZuoID8qvJeWb1IR/VWj3C8PHL7/LGpslgmJJx7TCtVCjm7yCmD9db5mghJJekEq+ATt
YSTQqDLuLecZ3fJxAUC+AwGn/oED2VfZz22b8ZI+YFx7bimxucxWa2D+X3qBMY/jxohaJEHBURUT
i8ZNolbXJi+m7ckE8aUPiU7SFpBJCZ9z9kn79kEVmTKwVUxtv/+dJDsQvS7Tb0Q56pmnjhwxCy8k
R+KHdGkzlQ+9CWt3nytWJZ5+mkImHcGEgk/BUWqB48e6K7cUSDHX5RbjeVZWyKC1/YJkpBiN0S20
UL1qo3bWH+8JDFmqAgD15sT+GYaPZGQBeX7IgPJpmmnrH4pmX3KdGMeJ+T20mi4EsWoDl1FbT20p
V6w5a2Y1R6msww2U8xx4AiKKfMn9wenuqkizq+E5XhW0fK14vfN2FIeY/JCzrpRmWPFRd9/D0aIZ
ouXI4nxLkt/W9DTvjGhbMfzK/Dqx99h76UvZen/vFvtrIkBVZNCw4NBJaXD2yM2eoKJEBXhgfk/R
2b6yVZ65QjGwmK6dNJKh7ZiTOivwLSZrtaGIriM8oFFnAxNqcrM7VRggCvLSxNXPTFCXlsCw72Gl
bOlyxJJdnNNYcwRdLvL+rAG4AoiuAN4aJBEJdj1znAwEErr/IjXlAl/9RRV+KMsT5vQgiQYyqj5R
3H8bANfRJbVHnhWRvQTGB9l1plVxTYuHP9t08zewuNcKhhIeFPheYhuQDGU1gehbUCcW4jfXXynI
F2Uf71t3nDWssXPYGJBY+I3l+3ut3dXgpemSUslBkcfijNRsNdgvdiJq+NViUhPXkpvfQBE4RJD4
ZQuoJQ2pck4lT99ZPwmT3EAz90WypwmTgMTRk6Y1yvGeEOm036nr58FBdXhWlaPRvT9N9SbXqirT
jk81s49bbaQrd3foj1TB+b8bZs5vE4D64039eMF13Pj0c7LmmbOoxPcKGFTr7Vzn23M1wLBY37Gt
u/BM2eov/5Y9IzxVfmnVoPY3GPNd3U/YEjuvdn37k74wJdw3gzsYPW5JSn+R/zgkBzuyd7RvZmzB
QwpyXfqC++eBQif0xomU2kmBvPC5ctAtyGAU19cl33tFODUnkRJKHXTkWaFpTSPInJ2qGHtlVFv2
2LI8QqG9+mFKJwUJLxANgATkTwRBF35RFZsra164fx/3cXGWrTe0SmKtvF3bl18Rk9MO/pdzZAgI
y4Qcax7Uh7txBHZIOs/MSb8RC2UCQGeiaSBSJQxzskSSO1cEBLhRfyPRj6mNwg/zhhi34cQOc5h0
6kZkn1/ZfWYg0GWPw1t09/1PnPrsbIkMLI1yRYvyI79N00z2cwpJ/23B5Paj/OnowQJAGZY3trW3
lrijyECmI1su6vjhy7TIA9pEkqy3S+LZUHVRJZpQZGQlyeTQB6yVWCmtdN6DqgY85pon++52RznG
jo4RC/WEB11WPeo9zsC3E65WmJbJxlLhc/Z4rz0dgqEyrXqEfNmMb6FKtiowpNDXmtgGai38QcRg
LfZr9FmqHnFBPTXK0F5cWFdlpeRsWtUu5zo2VySIv+vK+qKre2UXmqM+1C6gvrN/LJIhD43EAv2u
6moBpa5aA8XhOlKH6/X1nC12gcB0u0aIXU4lcZPMwKgf5o1uAzZ0aqgF4+qJW1i+seyj3R3V/JHr
j8wtrC0H9hlpwkw9JjkNoI/8/+FR2p1anZXCh33wOsrH3GtYRBpNMYe+qcr8MSynZ8jKwCZCMbF1
Lkiaisk2qKT1LV3J7pCCyjwR2HWQYOrqDDqh8SO4ZzqqzQh84zkVjAfSOoqjTHR9A5MUSjVyT/a9
LIP2Q0u1N699OoazlFnKn6qCphLFNTTEDMR0dlU4N+AK96F7iedu2mzwyM2Q5tIOdusJXcDoA+9w
7oHvlcm8dI8ly18SqBNd60XbD/Zq+ycANpDu1EnoeIEUz9RmJ0Vm69b86RpTPZ812GMDfTOpmoDj
gG42AuhJFDRnjOYjtnVc5aNjxcP8pwgekW2qjeJbAbQ7qzgdKbmZIwex/B/wPZjQU9QyAK2yYKDd
zp2CRa2wA3/xMCMy4G6qX6GOyZ0IbPsZletnlMvJslvbL5FEhr+ljSpckyQZ3KLrI9Fffn/Uyx7R
MRjM+xNGVfUeWnfTNrNtmSdVt44YkPwXCjiRxkxHwWM78+EERU0mByHK5mzY7C0ADuso2sQK6Iv/
LHCEvjAdJOHq+EiwHs/6V8We1ymr5+MzP3jvEDgMcB3MdNFfKR7OPUjG1l0Tc0Uw1FQTA4o1ssKJ
RWuzxOZuogzlsByekacx0xhdSCQytEq+4bgvpgrhFdWelUbcYzvkKQj4na9VE+X3u/ATSYf8+fgo
k6lJHkBEqHz+O8WNEFODIov+fQam6ekO/y33qdYQp/Lt2UI0ZM5loMO/NXpmQs8eozv4ILhVQsGN
UezLs/K0h5AF1ABT/QRVSdCNEO5UWSOTaN2iup64XHvCAyEXbjrKGba4dWCV4jelu/Mrd64B5ubD
Z6UJoNFJJ2t7Y1bT15hr/3zzaUwnC+3aSSFfWPB9RzVLodttR1MxFF0wKvpsFbDUdzcWbDRbkQfD
3Zfpu9OJuv2oziUDXk7sde49kHQnG6sN5POFYVrilK7Zlx+q86zxKTCRuQ1Gvi+qFJaNR+UsHvK5
loSXvHoCjAiCWNXNS4zCoU1fnOQRDzAQBMPs3SrcUOaPXIww2nHzfQymac/nOlLQAJMH8djjNME6
64yj2je4ZaGOLllQkh2gvZr4FQljK+nricoVZSpWM6u8WQdtY72d7Wt4wmukMxzLg0dvs0m+aolL
nVjNPDsxmAt0zSzSFxQ0tRAVNvLNupefxsSbd9WoPhH4lbRaatNWXJO3HTGP6tNhdA2QUFs6soRk
1khmwphyXFQ7CFfSQr0qQt5F+zZZQVuQI/QPlzz1oZJZPwVRuGCyjQR3gpU5gObvUMqWJn7Ad0K5
X2d8iALb/HlbsaPBHkqes8glozKjT1oa5pfGa758R0T3qTzzGTfXP/ViIKOfPMrY1XJmbVkrOGZ2
wz/uC8+QcUie87bHHi92mpXCMQL9zmqL30WRNgbSC28Fuy0mPXaSUT1+TM/VkaO2eATdDEJXLbr8
ECvVRf4y8kK1e+ZCxkOlpeVR6FFzSEc/5hh7QXW5dz4/LeLXJWkXcQBcOMuchCC7FwxpB4pnvjYJ
K43G/wksa8pf5lWe/+RaLGLz2qM0ExWVfFqKoxIrIp3u38gK/vYA/Tjn9nXReL05de34cF9g+t+2
DGc1tE3otNtgvz7QL+vA/K8oxJAqUFKM4CnOWp6+Mfa/6qpc7XtN7X3jAdkXS+GkJ6tjWH2D0hoE
Noc6IYdgRqR5xIJBvzAdL+W3h/OfovQ5clgpJ4Odm5eNraFxBG1ZnwTXfWlqH7dmr4sFvhCZVmNc
FZI4mVtucb+4jVMZvhygjDeYBr1eCL4orJR2OyFFiKMn8Q2ABOFsMd3Lbl4do5qeCpgKKxPEgdJ7
I4BVATYf7TxFz5bCeuAFxIGXkLWAEtq+1wC1pmViS8o8l34rwL4wMmwEvsXjaFyD5+QbBsHIeUan
Z+0Gh7I/ldgxnBkZGHe1AsIqnQFqd3VPSxbJoEzvCRzyogqKuRPK/gLo4xnVM4AE4JdrmY3N0r9y
sBnigWmTKqxON+82gQocfN85gLtQQSCVXyrXP4wuiRDcIH/6Bfikoir85mhi15nGTevfecNjBdmS
pa1MriAmnghj/UFrrRLTAo3teON2cr+FfFr3XqIxdzmbSaJg/2a58DYb9Mz7CAC7RQ8MCgsLtX6s
wMltQWrhD2/hnJx41505zH5LUVYX7C6Vxxes+ciDEKOyow406wPuNReBURcKGNFYKkVrHcb58tNP
zBGrBb/qYQAkySlsECpE8Yf9fy4AynTMTz6d4l+dUX+HY1ZvGY/ArksIlUUpdYAOnylhnIO6VfJT
s1ZY8uyrMzW8c4MjZCaNIErIc2QpSF/rDkzuwLZDMNZ88ePWTeBP44w6S2v+oBnCPmF1d2yPjpA5
tD87K7HTpNAUPQdsTqe96M9jrIgc9ByU6oA2u8ow9KvojN2kwLIhUDtokiKqHyILkwgiv/ieI8kF
PwDINrbT7hRWDLDl0VPQfMwmeU5y1CvMGde0UukzheiqcfGk3Gb9Ory41sGVeEvcGgrNnGzhIFHp
kNW1OM4tTuwZ0vyZ6yaR3VwkK+J+SZ+eIt+NERCWfHbLa4SYQAXInt+lByHri9cP0aPxFu6V3KOU
17N4bY0Vvop1b/29BNh7aITBClDgo5KnfjtfTpT/NBP2456p+u4p/DbJG30x6hQukCGECGVX0usV
SIdnd6m5E9JbKtyGu3bRRETtwhMj0W4od9yv2oUUZ6VtvlitJvegXSCFFq77VSe0+fCNQxc+Bu5A
MY4IWCcDqckb7pTaPJzWXs4lBcmpCg77FHBhfuZvLeUyB3axJQ2ZOfU1ODmEkjKCb8rE7qNqPlKV
IFN9t9JU7/+mdGbM9B2SwM0ZqK79x35/ERuiRgFDCtOLhapF3SBNU+wEscn6P6dkOW5t/32I8siU
3Sn++E6l1hDFasznF6FF+9wMIafHB4rw1EVkSbRliBtBCbvlJfgEhYQ6nxERBOZ2UFtd1KQRi9iw
6/ZIdidm93np5gNGK/3BzPipyoCFbH4rcIDd/HQQ31KCVfDJeFkJFfB80AHDBkAOJflxbrVKhCgg
4Zd6rZnP0iqmi5NpVxQZLXI6ESwuv3zmKRPbjgdDzu0AojMfwLgvkCza+LsE1wXcCW9uI7i5qw1F
XZi3jmvoDGZdHcxj3nleJVupYPIPuus9I9yOubXw8RvmJLDaD6cOfPecNzriajF55ICWlpTXYeZd
jveO4+Hc6xU2AqQeP5zQE0QnY7qX86ovmbugvWil2+v5Vq41YQZb/miFItw2Nj+oHve+tD9p2Kie
lFPVX3mAQGldDYS8c8XdyMl2ZnguHgBT7pwFjG+caS8acYVLRDy4uXcEyDBbpwHG+uefHiD3Lr0R
9jHPOQYkq+PvO0OgeKhmIfHiCYy8ykx5G+IfsjfMnRyGgA8i5Uv/5PZMok7UMruMkX1me+84x9dF
xWN09fRK1YfYN1APqsCHvFQpl2cjW6xmG2Bkkhp8woRMHQawUq6rvlh8TV0Db86CnJKK+tlmT/Rk
fkSYuM7qLs1Y7qyW4gVGG2L6RQILdB+nN6WhH4g4MRsvmf68ldP/KDJBhuKbGC1x9p9wyuZliywI
fBU1Bc7+x9l/qOao4jk5gzudSTHZg5sekUHTH3cvTieM8EgdDWuBrhiYTmi1muUm4MMILM4U/u9c
RStf0W73Ro7WAuL3sFS8FGKY+T8mu2KqBRl7o8wWVdl+yzRQkOHJmk8497M9wdeydnUzRyrXlG6H
VPWOTJnUdwA4HMjMc8v1ATJ1OI2sMQmOeO9DzF67584rpdGfOD7Z/cw4qK4JLDLLmsBUtDRq746x
+Elpvu7hmjMI0hrqPa55Vo9Mbhr/2bj2ePXNMunGj1KWayx3ORa8v+qqfHWOv1nj07NFoCG37C+f
fiGCWG8RZVczh98FiqF/01HqZ+Yxd+1JkeY+z8XNH2rkvUIScyw9F2QJGslL8ugxpoC0abL0NMPT
TOpcatVqVELAfStCX6ZBpBc07DWr/hcmnB3cclVj1IvZS6pRW/0R3C/8VOawTijEzYKFCWSY2mQ2
eiQDQp1e5PXTM2lkhYmPvXcgTiWqBHk/y15uUq1EzkzSFP7agkydSp0iPVeO+9NV31YHyEVrNv1/
5D8uevFP+LjpfD0Ohibm0Sccy2m+6xCRZd4BMNHVeSoEgiuEqJgsEKMBtk5B0yGgxD0AEyIJCF69
80+ygSexC3EYz7p6D1QXnEYANt7BsmxVO0ix7t/JgHGEhvGLUPBzOjITjMwz5QIQUcs+IYCOl0ij
tCaBY1ELCjvtl5XZQQhkMVYCC6E76xC0ivvxCsI6IUOEekMxpYYQWPnKXk8pgR8NvaQC6M12pyso
yGDZi5AveNBZ7QFLvkUf5qTl5O6MXJ8m3Onj7rBVrpNGUtE34sRKE/ZawrclQHk8Tu3XoqnrPN2n
3EoPkJZBRIGqVch0sS19OZ/wCB14dygQSResdhxTD+sJ6qjB99/EzJl1bb6bMGP4WTuXjmeHaDoh
KV/I+p96lA/3QUnWbDwUVhMFzOMOLcKPKeFWqrhchcwtVEy8BjwurZzs+vMyvA5wXfUDKmdpHROl
8HbJ8jOu55VjIprAxGro2DPiteKuAbiSaMaoExYPueedI3Zm1ST7jpynTeqPH+yIIgQCW5zLbPoh
OYLv4A1dAVdm57gwjgk7oLTbjtGyfF8x/pHies2EJcBN9FOlc1eZXTfC6bn3vX9jlRRbks5ppPlj
s9+2VY/lcpROHj8Qw510UhcknYQbSXksB3wcERgljNr+DUItcBGHDt28Uxkue7XjcaUHyh1Lu5er
dnFgiMAsSLor23Z/VAOFCLJf9d4eNV2SDg1MSE2R5DUlaMZrHeJgYEIzJz9ThZ5tj/MDWUxH5uop
16TcH27a98KawC1wOjniBs+Lvh+FFgbJ978A3lEYVgLge4yHTr1sRXTVKzaWJ1o+hZNkEb5S8k/K
iPyZ3dhmTb+NxeSoBXIoyxIe8KQTKVsMX91b+EisQRVQXiQDQKVEfK8XKNwOWMjF+HNtauPoY2pW
CW4jBzuAoo/+vJtAbZExCTNZ0Ywp+FwV7wYoBB28c2Yxv9qzGEjkbawo/+fRqtDUzzzG7+agWL9j
nREHQNAATmygAKqIlT81tzEkVeNNCqYqiGHEV9lCXj3gWGXdwyo8XJ4qeaZoTG1Byhv6LeNylMO2
EZO1G2VOVx8LKcU0HM3zhPDByY6Bms5iz+/jE+ABn/pWzfjaXyoTI9Awn2C2KE/7j/3B2un8ow3F
Qp09EPvfA0x9PfmtlA+9yU/NKSzTOGxF552tvoL9XI/dLbeaSmYu3uWgRsodP8GYfkAXI8gteKMj
gsxv12a033XH1749YwEVL88RYJLK/YWT9IITcSMh+EBVQibPJA1OWmDFu0xW4tnv27FI9hU6wrb/
ABDATPSWC3i2toVJQh7EoCFfAp0Nkc8wEiDYLgYHCNaKTry15yLmwn965tU67iMWDl1r/tlz0I8f
HF5CLKqI16mJy+72tUNcGI0wb+h6jqZZzFtyWLpaYGqp3oUjY5GwHiEcejx2vZFQK6GrTw6J2dMO
6j6w0II6bebxMG2pFTEjUWpV1Lc1A/VJ6LwpMMnToZIY3ituxQOJn06heiPMTxdrlOIT0mwH3nMu
BKtBFdlBF9kEmBoMBn8EatG++iONMHb71cwc2wKr/OYQLDLoRzqxUgeA3NXTW6oXJ/w3qK2xFgdz
U7SrQGRQpKSpYkMligY6AFfxHmEO6Z9/ySh2sCEwv/PH/rMZ3llEVAnLgQ5ePtvaInZAvNW3nMFP
L6/amMl4936/K49s3L57H0O6ZWKvSS2b6PrKFOMTupY+d4PErEzeoEc5g6j+euPWX/RpkO3/pDMc
PmXAQ7l5Z5KbAr/Q9f4YWFWiwTXEc0LlCnfeoMErfsAbMLFpfQf4tbi1k3FCHTYU9QvEiVsu66r2
ql+iG2v9XDzeUzBudq9x5LHCjHVy051MbJgZEOKUEpnAoc9leMc7lwDsNGNaT6euMtV+jOV9Z63G
YJspj8qwOhK4c/jwEOoehgKeJLZ2CSNJazsgJeKDGumI0pxiQ5l8p7Mz/+q5XGKUp/lM0qsNCyrW
BcRD0WHl/+POE9GbkD9QmacP9Igf8DuG9nKBf3K3AZNkPfitgi0wHD8JwXaAS+Br+VEX/XUkXAjJ
UXezpKJVgZbJppfw48CgtHye/U2kd1vM8Eo6WDlU4BFIuw4NcB8sST1g+OtNxTWnD+/NO3qMPN8r
ur0R6HkHSux0oE/Aa0Df1H3XXkqALwd3AROn+1+xlbrs1KXvYJztv2PyQiiR7Magvd1G1JfEb2wx
EvjJZwxF/wsCHwklIwHxG4mcU3tGCB5nVkP6Mf1p75ydhV4PO77wXB7tAAagQvMVTM0EQRkYpYwr
/qT6LECa9KfHB/cXg0n/NVpvMRWvE0C7Wa0Jmm+E7GUi4J6OfUXqDnzz+YZL5QvIr5jpgHYtgVcN
9YPWXDmHj66m96m7buhqUGHFq6E2Ul83UXLYtUm/GTuTA1ZsI8gwdgp3I/qjBncocU7DDz7t05rJ
VYC01P5mQGYx+BuoDVbL5bF7jHyX8/UMB3G3r4nMVBFvzVrRfXFg+0h+zk7r5J4tSOXTn7YUT1Fd
yDhS3nWZL64N1DC78OnV40pKEwEMuRIKjdSVRU0/BLsQjIN+cdPQdn2feFJBhiioDZu+/yrLxyvX
35COJYmAatvnrtUXA7/jKXNOE4AxEK0agXLilnXqo8VCY8oMF4HnZ9seiZOph7Oo+5ns+POpy829
T1Q/LZ5aDPlfNxuQX6iqXkt9tJdZ4kCf2nKpfidJm67pxlJaLKroTivbbUnxvtUyY0r2el+EBRHT
rsdrGLPjzuzysyxPfSI4zJZfk41DzNJvRyWfgrj1p3VWljqfEEuOxb0tcr52hRtEx5mpcWsh7M8M
mKyyyET4H/A6wIUZ0+A60XhJeewjDDCke5hyBCodS7a96+QtqnYfZ6LnrNfrxiWCxt/rhnkWzGPg
XeAiqowx7fx9OHkmbg0ibk1DSkgPrKzovfPdMNqfZlEMgeOfgEFe2935veeZGN+A3vaU3I0n1BdE
xCSuAxVnvyMYD5yFzhhtX2gydDi3LV2sWn3/9LuLkW+E19JIgNk5rtkyW+YoQbQbtPMYToFgoKOk
5oz7MhVjiOoadNv46dr3mELRORh+OPX5h6mgGQaE/LgQp4vMWeRixFq8Qpwe/iClZbrzgfGvCfRe
2cSV/4gARod8NGdwVLVPkzvOo+k50pM/E/8xoILe1+PsYw2VKs6uYTP5szqR0Q5eG/jQreWmrrOj
Gl4Kq0T1Wv5E0t8YSMVLSiKp/rC9UcmRk9XXc4bPRoDGh27EUrDPGQTA5elmw60C/YuhH0IDK33p
UdXJVr9JZPI2pm0KwGetNTRi/GacMZCr/9SbPk9YTTA4GnUZolr3KRd86wSRVqwPq0TOD356LX+J
7P8zJ3L9ZY7Kt7gusL+gULDrc49+xlyIEuyaWeIlOZnIKvI297jVogm9uEe0V8lM+tGhn8GWzuNg
mlPIfAVtWeOnxB+XmX0bnUTNYGXVqlCy0ZCCML7fSNWVHzyTqqYFezMFVdMgZ5WNN7CgCUGvJn0g
xEKGgGI5ffllqmAYmW++N5AARzKkPnwsOkQvsJEkpwlTdP7C0MUGJw2FW0AOPaUfNjrNECsMvsQR
KRJi+175ZNwRLVFKmzSvBGZ/UG1juetYyF5y8JCkZIw2FvvrHpOg06GpUZBGhV33z5sH/eYysqiB
3iS444ec96uyedRytyUIyII7yS7kahBPlCOz6h4O3T5g3+uWJdT0hLIklD5d4r+SQmStgum6/A5m
KYf9CXi2w+aKC90Psu4sST1XlrB0hIZkCdApGB67cbH3A2xvkGISyNd4dM6VcK86HfaKO6GHj49/
Dvo81R5Q44vsdAurzxn+23VEa5qcb8D3c3W5lvdEJSCV2S0NspO6pYe4dJ7LTOSH21U4CrEvLJDp
6haH/b/yX3++6Zbnv8AZiGkunnZc37uvkHeST3G5CfYHgw/Qzw/JpUESRaPG32t6zMRKa5pFCqx/
UbJf6jy43OUHuLoU+ST9izOOgEIzX/Te3ZmXnuZZFNXtSvupYR3X3x8zi8k1kHodafX0f9Xxapua
FJUJhKctmJSyxoikVYMO5LvF3fIafB9ZgWxMs2xv86+eFBTEWqtrZUxF62l4Xf6wj5TlMKYsUZNx
UIg3nCS2pwPrrqeyWkTA05qpZzyh4pub85b76ePHxXBVEmhqnDL/CXIE+kUWGBY9F49CsVnnvG93
i9+oF6zE7IJfP+CTIo9EOOWztItNIFOh+Hled8fuEKLJNUU9/zTZCoc0mcgd00JZIsB7Ta7buupz
9SjWzDfiYxXNI7+GeIPK3ELUx7IOUBNarSNdQUhD/KhuT8DTmPWwdn7aVWxaWAnEsJblVxshm7xz
mjabim7RylBslu0s9/zYqp3E/pSEqefxFgOKfhVtTAyCa1s9yydIkvsP/p2EeMsz2dHmXgaLGqL5
N2C2x7PND25IKuvJuxHo8sHea6kKqAtLKMjs30gJRWIJu1lwiEXyZIYAO2Z6R5YEHIdXkrn2bQGp
HUVTCNECCp6thkLBkAL0IRhfIk2ZkKj7iJFcIPtd8izn0qXrOZsr9sQIVLff/gsIgBImiLqyjfAq
fXG9tniBYmf00/VxK4NI0RzUfJw9Vut7bm2cSZJgdFu99Yo2EdDHongvdo6LHc8LkKGbI3yS3tda
/8MxptkGYLd0cDoCANbcSa8AKkgeek1RECJ+9YsAk8rMUuLNJLr3GD6LizohoV4IrytUN9lBRsLY
DEvXQjPdimjPxS8sY0+xbsK8pjvzNw4UAn5dWjtO5bNO2uDDWgejDFXBccB9z3fbclb/seeUyfuk
FN/i3RHA+Bo00/5HvU36S+FTmgx6hHeJOxQaqtk9y27SCp0QC46N+K4kBlBIx+CSGp0rVeyrj3Cz
vA814TVXFSgfKWjwnALxJxQ92K6TCqH4lQjfyfVDzV9FeMqz9cXnLXT1V+eCBORAWvykvzDNHKyd
EZnFEB0h7PadX8cZOm5dGOx1SSRmcPW83aRf6dee2EhioQW35bwX6xhnougt8+7JacMOJrbEgdlQ
SU2nIXvrQ4u2CFVI4O9iIVJ0LBJAnlohQgFl2sdlpE513XU/ZnvSy+4xgrfbWCTVdEBPpKgs/zmw
jlpuMA7YdMKQku3omx3RfgCpE5Ct0gDZn7iXXIox86CZdIfFDsvLk3XBNo+V+eg34VZGw/e9ISSU
BWwCuMgFdZ3V5/quZdgyL4HBfjsLekI9iDrC3ZFUn76hqSSQ0gQ0bidlnrgvSPnw3itnfUyZWq+p
TapbnX5kfOvr/Vy3Pe5jesQPhmWMgWSOXJDmfju4cDU0NXl3brHPC6p/+0wC3H8CXgmCHOZ/n7a+
rdYhz5sudHHZwaw39NCYHmA5AgQaeN2P/2G6OejDgtv/82qZr2o98ApbeBVjYtJqvVGp1aCCdRCf
H92fMJzxx+Ei7m9LmwyylpciviqtnVxs8v/VdwhcWzuxl4F6FL15G2a58PKp1iMyjgBPpDt1zurv
dxa4iIsxhb3b0oTCLu8HcIOtP/dx0pYcRJBkJufwslesqFRJJUYxQWrf+KGQMWxVIO/Q/qf1yzvP
AXrpe+faMQvdANsQgKX50Cw7MDEigFGvrIbB6wJ3KtFe2hhmidVhgkb0tw9CZfPNrrdZE6QqNTEI
Ao4oBIA3vps927O39g707qSv+llrzLAeb6Ttizd/Kxyh7AVUNnX2wvLpFHE7vXj3qh8psjIYEEnb
4xdP7JiPtz+o7gJwaKHD/wyXNdlVYDUaa/Y71FVfuf19nAD6lglSkcGdDcPLON/Hxf1VLZHrsjHq
5+dNBTIsMWqvkLz4NJAvcMpZQWVe2j0lKkSWteCEqB1fnaQUMNyyUFtS42BKuAWdbFzeOekWzGW4
2OqER1Mqi3hMeLHFzH3naq5S4uZdTdY9IOmBWZHTJ1WypuRxjMs8pRqgfar1lcmY7D6A6FnDwBKI
jsHzL48Uf7zG4HBpezcP5dxry1A/oN6p2P/loKRqh5zXri2fAAGAWjPSIOrTX/Ri+c2ebnfhcRPO
frfeIL4JBhhZ/Ppq8Oo98OrR3fSFC/7FW6mIF77vMF+vYWx3sYxjlfeEZQqBDA6/WSXtQem+s3Ff
iB1mfWIA+JK5F8hWI6UPIZxLLcnv5c6smPZ1b9Y47NjgBMsbMm+HcGxFeEZ3K54fJK2EAk/GqtIq
gBieWrsHZjLaspcwr1rhdVcuFhAluNkehRZLo5PbN3mlqGC1qOgrnM84G7Ixi5Qg3iZDZc530GP0
u1oozRWSSZvo91miw+9hlbMUO9qhr9nTvWkDUI4KqAqOghHk81tyf5xAEzw9aybdFdGpBjyn9T8g
gPvROoJrkvwiD/MeNGVqzpkYTzU//8ynTuJWixSvRG2gw+yhV6kryU4+xGPwGr3/wVdqfxTHwXuI
CgCRPDMAHCGhFs+sQTAskLl7NjYhYWlXZt+2vA8JYw+Jt5WyolTJ5nVm0oizcWj/oIfi8A72pz7b
UHwnlIT57I8tJUbiV+d9uGvE+FipZreQEVq+WsHDHU8UdoS6CBEurxfSMskI9zNJw1E1qut5FUW+
oiy9hN424v6XGRoASpQboc24ZPw6Iw1GKVL9QULp0AyG0DPBDrIkiGvICKLP5xlXvsEDuY3KHJf2
HVY3uzL3f84n1fAgVpOrY1+QPiCuFM9WdwqM7M53AdOrawGWNwLSEnFXObSAqLqi5fFt72DFAcaI
OcuLSyMktNolGuNJMcTeYALzEX5PpcJuBa7vPyDscf3bggvMweCTQPuSIP6Fhmw24Wg10LC5gSbV
q5hUrII76rEK2r/3jh+H83OoVEmRp7xMIBHFA88wpMXO1NiUR4alJD9IAlDAK/AkD+eU3AoOYuaC
LDgDTnT+IXcC7CUiMYTZYSP7Q4pdjEVEmmC3YCsIrdAnE4KrAik9D4CExVcudnj5z+ik6p5oxP0B
w6jHV7ITjYHNwvVeZTQUfK+oUSPk/02037Fh0UDmTBAq2VlOcKjxKKxU/S1YHKelPdUyfI5txSSU
pof2USSBWvxUUsdaAExCC6qvtbc50rdYF/R8GMAhNKMdvmeJjXeeHjAlF5ndTz5QkBAr5UYLjcQR
olIES4sxHb5tb8/3MWkI6VSx+jxQEN5pssQuHCAKi13lZo2vJNEzJidQsQhvAA+QbieMGQ303jLl
VdQ7Lq1RtnIM1VVCmfHxKFCt4fe2xpi6buBr4ffQjY4aMzchUgt+eJ3iHTsI9Td5O9Seyni18Fit
RINnuqy7j69LnrL9bVmDoaL6Qku0ojkmVCG7UOssJq4m+8UyHb50GtnRybR8ZAULcQBpLZ8BFWba
lf+MbiNUZXtNlVeAOyoXDuaooxgy1xC/e4rcHGr0ej9jQSFhaOTrepAni/7OZWeINeubHpHRU4X6
HaYI4v6n1rPeB+tSpVuHn7hn/JO2R/OnZepQ+NwKQEWyGOnvYYR+ti9xkQLn0nkFOLSWB1sYOGcR
ow11WEKKNMIcB8vo1CPi7mhfcUdLgSqerGPJSLZ3MsPBmsP8VVJR2xuuMWWfb8khx7fbrmsEkgru
XqYdY/hWs+gVhURsZDM5T/7Un4Ejrf7oLIfT6oMLlwu1pTAda2EPorc7xVnu475FhJj8DLhL/DBx
KPRxdA6CHd2WA2G5S3G39tXuFELxyNRCe3xu4WNjCnBj97x3dFcjJOUv9oNSmnA93DrCFY+AN/iT
zlsr1kTi2l/juMlBPaIEoxMH/uwXT0K4lIAc9aDQwDx0Js8UDAj3dvyscxzvay9G5Y5znkUsjk3O
lQl65VmtP6yoTTwMOLnBsBIFrg2Y3yB7BFzk2uMITHoeJOWqR756ytv7flRvDthIxVaGIkE4g4h8
Bawp3r06//HBVWeFVOoWI8IEsKH7vqX7SF5lsBsYNxRVW2e54cy8nux/EIfD6htASTYlh+JpNhJt
pO8VT9ukejHix0WBqf39XJMHCocsaK4vHLykxrotGLzEs+HTf71eZjekIeLNAtXzFJsjDsWWUOGn
ixpBvSWE4BDVpo/uAPzc16RdExXW/4+/ENxpzezO2WebS3ffsa+OAcPbn7iI3XfTaxMLJafy8USb
U9dvgTzRoZCvFN6Z6iKPErmkzQb+TCrS/jj889paaQCzN7togwVcXW5B63MQkyXU8pENxqmZPWxG
CFQzKA2WwCTHM4bcri0Zky9q/Kok86pSAISAyQOQ064sJUUp4pryUmPB4iGqQB/Yt+bXpeoX+9+C
5EM13htIa7iMNQL/yJWih7OkoKcYgh7wrAW2Eq+I4GHhu1jT9KnI3qAfBAjNEUe7WzoHd9bUoh2O
c2WyrTAuqBUWkBBw1okdwqPllBDcbuWF+6Fcdyyx6gV5MYtVHpSHyRw9RxBNSliZUGXDF2F0DIhb
9+1WltGWiWn2dvxtY7LiZmvomuLTzcSX1/b/Ugx/uq/h6xW7BqiETaUGdCsKU7h+L/NqO+EiG17+
6p/sO10KBYNHCxz2aqwr9s0yY3g/Hmp2FSv4DMXpn81DHXPPbsatNG22XJ4lmFH+gVRkumbBPY0q
m+t6b3I7xCHeHhdt9ihf2JexBMGB7udmm54Xd9eMR500/p25knxKiEU81YF4afv3Vg8GJKtOCGSu
pBzTHtC07WMgr/FF4w0PR1kyPAM9ymSpbimNlX36NzYunmK4A79qS2Qk8hnTqaslXlBlp4Y4VTtO
Xxj84DMHbuppxylyQnhTmm78IVxzN8VWl53PxHSpQK7CQp1FQxYtDY7VZWRGnevc8GlHHDR/N3jA
O+ZGmQHEfysdX5/DOG0+w/qkXDtjyygunLstUKPB9rn26mzXT3Mb+7DWafi8HKf2cT39D5whI/xm
p7LlgjUqojbgdM3c6X6E/1IpNmSRWQ9r+0KfxWoHLBlwm/1ogrW4PWIvaLUjj/jE8+1Dq3j2nsI0
+qaBBcA8jn+XpnbVS0Hknob88PGDFTkIUObrjo/I+/maXnypYWwAIFlJGAki3cX9cbc8rSAGA+Ao
qxLZq9w8CS73/RKuImb/ikd8KAF+UoS07D8fVxbgXsUczEZeTe86uniCpRrzPvpjsTCFVaBa25qK
qKBl75caPzBa4sG1H2gXTwUXnYDxkqODFe7nADwyhup/o1rF1slVClCSDu51nlp50OcMi074kMXO
OUGetLifeq70C997kkvvEZZ4a4cE+ZFRHEYNDva/F5k4bMCxUjIrrsTWaWaE+Wrgv5xABkTLkMOP
9oET6q+Mp2AnLn3QlVY+TX11Nz5v+BWrF3WzIQHYb4ckCFCGfbYujeZqyfNNREalmYSaLysGKZQa
amNeKcxa95/W0A7YiC66ZHQ0UXD+Mg+uBdmvNGuO11+GMLGfAYiMMU7d9VmjXkDv77udMNb24lIr
aYk0VP5gqa3fCv+TTkhlAsQrSmNqBs3Ra+iooA4nmnpqzC0DoQ7WaI3Khn9cURNWMS9YW4603Ztk
2ZO66/wiDFSio+gAQju5OTx5okLlkT2skg81ZhdQclEoSB2Wua9pJKLqSS8SHX+C9KIklRRNGZDQ
pMkVsxVhzjr8YHkmEShmNekdJlftMZkvCSCmGlgKReEGCuS8wRN+ZahOrUhPJCKLPiY7alIvEgRk
Oz9/h+XQrfKf4ISLZx0h8aXRkDx41RNZsl/kf7bnAvhoc6/scQp/Sbz0a3G80bbnwYhjTbbU3phq
EGltliM4clNO9e2W7DYQpcEnhg8zK0P9VDntmV7COvYZQc+QublyNpD08uH1/UmxaXjMrKvg4NGl
C2PG9xlqHWL9n9msJICJcNFzc9KV3e3zZ+79mW8jEnuWlPH17/ZqncIrQG6xzr13oJFBw59aQyGe
QE4zxiGUyOsyQDb6F/Co1D45DuwQYF+fpbQfO1hjvYwbbGyuaNOxRRQCnfYIgOYv2j+jyGGCVRfh
UZsheSm9m+bKvwJoWW3mp49c+8kbdkYrglXHgXLO/f7oFkRrIwZM1NXuhkOyH3CMKHU8itk/htXX
805oOQ93dN6fDWMp1DVz49rvBVtmTPwsi/SSfO4LO21pS7RA8lcFFVNAMN1mZx8dyfpM7IPFz7LH
3YGOdknKVT6CbiB3Fei4PD/joGQTeuruWp0FruXycx2K8mFPGuctYRkJiYjJkUDNpgDJtWjIgzMz
jVTWws79Pwdbil7IdH3/YL0rjL0AugEJgOq/6CJUZ+wqPYAnZNeKPsHNLO7B9aVf8/T8QPhVd9Am
D/cbHyBSksrjy30OCzbPuG9O4GTOsp81RdJ/ogA0vBu3KZp+VqRYghDJ2LeuGKkAOJmhEBzIYK0x
ke7vqCZn132GJt+o+bSfET94pxGhspAzLOExXb/si6X473so8VOF9GkXySdEHOE3jMbLqAdl9uGW
CsZZCa8RGQLn4AUPEqPZyzwPaf3WV4/bzGl0Hs6fi/0Xrv6hs1r4MTaEs/ngV+L+qJhQxADDLksH
7xwY4pZzyN8+DbSnWvn1zTpDQ7rX5eQZEuWqMTtnG6zzd9oo6fBopILjBvOukApxvN+nqmu02Pis
RnIvdaoppddd9mRUH1qUS8CyKWr+vILmWX68vNrb03Rd6iLZI5oweKRR9THE8zhpt2TgFCopU1yD
uGweQJggLCtuWwXQRkQwp7vKm/JXyidV7E+l57rJuOvVK07YuRTkwNu7G6AbhZAgUNM8CLkti6iI
yBR6ypigbBRkZ7+i44Xsp5G46aD1SoMhUdd+7OUzAzMWe/D3d+KgEpACiGcs9vcZwgoJOhXNreyt
Fyrc55a9pI7tRQM0hoq56yPi+js2n2dHSTfEAj9G7stg90wDENmhc4DH1L+GbfLPsUvKTDdk0G25
wRCjBYuC5F4VAf68qebz5lHKkpXDcUIQO+BHFEaK02KKmzexMRdXPLC7JMeJR3Byk/B4DPG0hE6B
LhaUxXrwZaCows9jlWqxfRtk48CeLUn0wgStPS9ETiAN4zI3kq2UXdqGUjjlYLlm+eU/z6GHf5G2
0kVJWUi5lZLtIHZN9FWabWPPlss8OUr81BvD8DXpuTOvtoRym3pCglhoVQnK1cLzlUbYvQbMYlUf
xRqedqyJFEykxgsUN0qJgUMRviy6oXTjTPlOWDbCViWb0tYdN4xV1WBqdifMUejNrrKldQ8wqDln
5hmv9sYC+1AlUXPJPD0d/D4JZtdYVm5n6jPTDzodUOZo1t6Wk6ub7yAEy53LVciJb6ZZILWZnUMY
T+C4xkmgY1HmfgAsWVtKXeOblhXpskKKdBEJasHd4s6MkMzBEukMeps/m1OZHr1w8IPzZ/cA+MfF
uWuHeTSS85pqwHmgtHsbpicoZ1La8z6frJYIaDAjiUb8xleZSVREj7SupOzvHWS7jrnLu0QF53QX
rZPHzDmJyJz4bb5y3CDxsrP5hXgoGvB+L3LRyFiTET0CvAzrwAqAurXoa09Mp0o4hcrCBbqgxUk7
ZZRjTxpnntVzYy9M1dMR+ePU5EP+YFdjpME/ocel+5d4pCvYR0qdW7mvyCOV2MH8Fe0lhTYceJa5
DwSqBF33D2CbxRPKADGr77n9TfTi7u0sdmM9kdR2pe/NrlXQPzcyzB7tBh0maVlLfAg+41cWVfGz
mEogG79XIVW/jcNloYSpsjnlDo/zwD7VuIbqmy2F0nq3csAVuxkG9UouWx2fWi6Cj7UHmCLNWOtj
KonJPUzekl7ii5JN9q0cE3XhbFuPh0O8FxjUjAX05Z8hqY8b7s3evnvtX6ekFSjh9TRqMoosAAbN
xDQe3cOwNFB4fts/goTXFr120Ynf7Ygs1L/Nu1A4A2qPoRie1tT/+CAht0jsexFhLu342gAdAzjp
wjN0uee2BqKIeMhnxMTvevG4YQ4yaRHb6rWCGlBDnWsB5oqlZWyOv6wd7iCMIyHGfSFiKkFZJbnp
iI4S85x3P/CaKSoLbl8hwRGndaFmLd8RCmyqrTHsToqoYfoXgWNBaaQ7XGkah7EgoJ9tvPZkxYDA
7eEBQmIkx80z4f1Def1GC4hltSjH2FqKRHkmmA4VBlZyDepvoSXdFWBxTTEeCboduHz9Oirel+Vm
91WkZwSNERYRo0sIIzwAyEXGY0xFs4JwlnfmOEOwgYwpnlkrhnO0hZrsQcleUG/QdaWhy1bMH07x
IohJzSGgORBHNmDXudZslrd0Zi3awDqcgs8TEsquLgDJM1yNVWcHNBxZ+jD3TgloJPCJ/9GefdJ3
fRiyd3aN7ZcRiEWjz2BqDRFzuSPftx8i/1lYHPyzBj/r/MZTFOTz0vNmWS5zkQAATIJCwfS2xZ7j
RI8sPgtYMXXN03URgcbwjP3o1LCAQKDPuVmIDVT6JN9P8l7AEjQ/2rBHEp+i1RbJOLvZXCam84Ko
iZ631oTrIDstzqIoPY1WnTDQOoM9kfY3oTsLETPVAxVta8c8PDASF/Be5Y1QNrYKNq+OMk7ek4RC
ktCQj6sRMy8umAJhvQOG9KICT6QvDZZF85qtgFSTLR9VB5HzgKeSjigshm6ctIboeRd/4EQvAVn/
N+qbPUBzYRy5mEV+zphVt6WwmOdODZRvdhtMDfDIMbbGre1f83j1Tbr5/K58MXyx+tIGjkJaNyOZ
dei3D+wGXZk9lpvL+AQ/cQaT3yLQfuTtcV0Ij9rE4bTwlNBEl7n4OFmxioLIyg5CMx5BIkY/ReMD
vnOXfL/imAy70FYKF+YoPyqKQQPEmu6I2getJTJLHeeuqeobSULpDXq8ze668bnhG7fwBp5BDG+n
tDhYfe1JhEpQ5vDdof5pDMVYDBMH4jErn1o6lbZ+WtFBXSPp9lpf2mN3q8O1f0W8yBtkgpkGN9Sv
FnbFc648pohCQL/Puj0ID+Vr/Zo58oHRd5MdjfYk0GcNdYke3QXyUZg+dXct+pEzSg27C7Em54rP
umhtFiQWDJamvsK1JCuefvkNG+/dfRPQwbziWczH8B/5VkGOVjBM1kxzff861fz9pkQIwBVVHOie
GwZHMIeC/tUrUId70FxqQ54P+aOb+8iDOFnj03dxEkVv4Ti4gmNse9+yhQ7jBvZoFyJND1CTAZ+3
9lYB7cbgNk/Kzku+mLcMNipfhPPGxGDIDP9TsL6qPoo3rro3z5jQRj8YCjWBEUQ7QA1whfKTGs9i
l36urxvSTDhE7zrFGK74fivcWJkOcAMwhapx8gkp2F1HUcnMroxOd/3xLd4OclWhWQJWvAFnU6yq
xkSl3lj/A8XsQsHTtow6GMNLNL6MAJyVsU7dq+n6rfV4wgqclzMA8OfqiyDbpSXZ5hceYqaKzdHg
cPupiff5RL/u28AoKird64pc7+3MqNEwQLcHtv+RbgwwwwF0dbKu373RLhiCtwsFuKEAao7ip6Gf
TGNr5ktxWUiZSC1Yj4icMGCODQ0zsP7w5zre/IlTBhkprQUDEr8BWuPGFrBvP1GZrCtG7lW9MSVe
cc42jSH4oC9qf0Fw5Yw5i81wEhAGkxISn9Lh8wTKbFG+IA+RysmlpUUxNoCyCwWrRAg79yNJ7Cl1
j1tyNxaLvIyeqoLuf3kd4Auux6RPrl6WKQOfK6IKcbkIAI4ZI5cRWQed06+FRI2WZCmAIkLCWvTv
OOXjVfKYZ4ZTU3NW5/55es5M/45C67JXXQ2ogxDLJeMt2OZdC0nN8VnPWQGqKM6onG0SG7rIaf+k
BxcQ2VTy16zTEcQutYHJc2/kUKdbTFhdTRxlil0Drsu+ZtiCdF6P5zSa6PczzkmEv7L5HDCVKqmV
1h6aKDds+xXBwtIg+CmIFXhJsxma4EbH4FF6p1PnV7kOmYj5gb9caIirE/FMyGczkEny+dDYiKUQ
RIqu0r8Bu/irbBixcCFGg+RUpNOAKqx0S6cHCmIQpA6R3MDHm2T3UAdW3olIIi70Vsz0R56UoJHk
2kOjdbcntxSyMmuQSnGe8ePipysjLBckwNVbjzvFl3giS4uaXpzM3Wd2l209WdvYWBgkPo9ah5Er
06jN/fbRW7SROpYHlsf//bhojb3oAw2eA247Yv/kTKPpmwrZhIfOfXEfkPXogs+L9bxztwNovRVp
+19mkFNu2gCustptFBcRPBU0C7X/eZG59DZjISXLsFDpKJTH2O3dULRTKdrqxXDNx3SqNzEfY4vG
6551OanG5GjZwC5LbRqwwe08kyhGSWucxGFomHXYP3iwLc3iKqhn0df4bgScxe58DnVaY8H8ayEn
8epB21jKm/GDZ0vokdraQi1Hr4NokbnTz8+TEZwsSPewrv6mmIfBB2hoYmKAnTIr/uUm4cjB/zF7
HZ4vJJqNEUniH7prRUxA3cXJxv6FSXyHbKiQ1z8qgqF3gzPy7yUFbzRvj9NnXENFFEJzAbaLB0KT
lrxaS8rMw2KP1cXXgTkD05daqkwpexBNRoHofGQM8tVgCRCXLJTr3wE67r6JnkzuDg9LVrw0XaOK
trGXLBatxIHmbCDA4bCJydsftUCwkuP5FglY6tMHAAwKJfRznk5xRahywoZxxCeKF3xy5j3xdNG7
GAtkw6kK8r3qSiYQY02TUoNMnsjTV+nO4RWQUf83rp+ONLkSjlEoECT1h/nt1DVfrHOYM/Lbu43X
UmeEDfWJcdQM2n2QcdUNkgzozlTrgYsMSDfEGrL1epAamqdqQlf0qlzBah6bdbueaT6IO3WFzyQ/
93zZUyXlvH1G3Ti7B4IaQspTXnnjnjWRtbFQHf8672TUksjMl7awc4pIKRG3A9xlop5Wf8qWJgW/
zddOofKUwoax7+Ar4rkuMCyCokCWc+xqcSI3hMlRJOAp/O2CmIcsD0KJEeodFP9Tl24NZNYFZWpT
zeCVcXnlLa9jfB8qZ3yrPdbrzKE1yLV+XN9/3FrcG2FpqGpEvf6EbO9mJYtUdlbaUEPs2ST+AXsl
mtkp+FQl/pxNaBZrXVdBz7Ix9/Ah4Xf4zohswigZXhCbLxln6eQU0tGdrWLBnM+6TPms8XSDV4in
pxI8jJSyeKZPotehe7XN1RFqOhaAyzxI55fsEwDPmKNNzqNQNDcdpZ99h+z4KH5NM/AAAqnzOMSL
ytVkbYJJkgZ5idbxyfdhBTcWp6IOqgxQAp+Ax8pziU4HYllRJ5a2zXcXcV4BscaLX/iVpo7Wsjfj
jDV6qe5BuNoQPjXMtTutmrjIp2d8iuPvWuw4f6XBSvRM543tKuHaAmzgDjgpdtEMkJ/0bGbf34+a
DGni6qk9trkZc0qZlWfpO7IEUlxJcex4Sa//wkqhMNbgdEVlOGdEzTywlLe1zcVlCeX2KtZsqhWc
UDOtyw83nm8/kNPwKqitaAR2qVqq1BdaGhtx1BzMpcwzpR9idLYP+FbVqGgnMeXvCGEe+F+9s6et
EraFgYaf5mhxndgBbWbBwosmIPy4w97Cb3Faqh7Od5+X9L3rimbGSCZhGjh3fuNFBWVjAIz+RR0X
j5pJJ99tBArMGZ5riTcDEMd/yIzIc9qAMBIGhUchdiWfVe5W781/IyaTIjbK/ulalJx1TZ37MSMp
sKLnFnB5zO9lxWuO9S5UUi4ddAN9bFd5B+smcLDdy4W6RfyyOC/GjhmxaF9ZZkKBU5YJs1iim5Xv
veG8CLJudQsMy3FBU/E7/7b/XrHcekD06WCr98UWShdEUln4zP+DdeEqC2UnLRW5RX2x/lusGKwT
aZ4PLXqgDdeb2NC8zL8LwG5Vdq8YeNevxavfSQD2XF7jAyawjMJb1F2RBy+W03CRYC+LVwMw2n7E
RzW+RPTTMESziStp1ZmBgTK3y8wJ8FUPiCSCUDnJ7zeMnxxXZykUdgLhhiKhgnST59P90Hg/uhII
Eup5IrLnLngzj3pFFS2shKel5Q56sfYlllJ52QRtYrmWGbtz4TXEJKofwaH08BA3acDfWpVhKfaq
GlfMliez0GPakxeqlPbxAcQJO1e0MfwWout6c14DHQO+JX4w7L6yP19aWQ6YxJ6Irzf/SboBYcnK
Um3yAAwTn1tO0Hu0c2T98WYef8m8qHXpBVB1XPzA307Yd6sbLsZg9KA/Xcrtkc0oIylZQDDd6YNr
FU/fQc50sBdYgsUaS4DqEg9dQiBvgEVdUytpWH7GN/wie327DR/a7t5YhaMikg7MdY+AxowUFdUI
osxctoWDfIfhaN5jdkWZel1O10BM7N2MR3kzL8WdoUfhiWjDL+awjYY0a+cqG/TxhAdgbxkAJRQO
wpYloNJR6YRyesydlVHw+X0cIvMx7BBtABzxAnaE9IRUlCrou9tgkPheFyrf/voKmxpYXBdXL7NP
L24Oaido57qVJxbeakruDutCpVqT2Td8oDq1FCGd4cNn3Iqg17UIusU4+hBkS1NK5jiuRPp0BzO2
Mt7BMgWqfufOBr+bJZ5XZsMlDyl9IWItGu+JMJOomxBkScdvJ5aPXK1LMI5D06tlW0a1+XsJkoxg
GAOgWcxs2HVTZ30Y80VjxA5rVCsH+kcFI1lCtk1FAF6/Kq81wcvOBJWtO+NTUUzdmEwChuxHFfEA
teg0agplZ65iNurXOPQKv29T88P34FaCBQz1McqLw52yHsyRUgSzwn1PbGwToGJ1Q5P/xyjmYqN7
jElR48++tBXx6se4B1RacSuLen+PxgOFqd7SeaKw193TPEvv7JUWEp28386LWN3ypwFzCn2LSxWV
uYqw8JuxY/E5BKxVSuQ/rh2wieyu0hw/yycYghGtKc83f0wphthPs4hBzxifyKl52vhEOXWxpse1
pu3i1t+PT4NAPRhvZx9uYM8RidDkz0jF85JXF/NxZAELGe1QZyvG7bTImRG7s9le+OgVPYyUn1LI
cPKgSXqEXD5ZWCI8CoIXrX2PpeuNUX7Z6L2N6TrtuobL727qKsJieRH4IL+03L1Pu4Fd25G3P5Ck
Ve+HZ0QIkRhojcCpXKxjCWUhPvnGNOxkoT3P+9e6+ybIW1F+D0JTf/ySSjSU142twvKIr6XSg5l5
6/korpvj8Yqz6zZ+rEjoT7aaZ+0ZBmyL9hdqLg2ioRpN1B7Oztm/CjQOpfll7tb6MiC3TDWGGySi
W0WNBbh31OwJE7qIyee/d42iVwJoVW6ureRUJzqdyAYLoFc3oP0hqdfqOg2rsLXkEOZyyvmG+gNa
RwLX4XZrRSPT5tsAwKkTvrV1VvVfGiKdgm6qYTTo9EN6z6lre5WjXlzKIE6eoK5jyS8jI+hMywnp
DzVD9HG1Y6c/l8a7dGCaz6MD5lL6tWbMuWQJd5bE31+V/+iXUh2JD4F9/Ea/14srFhZZ95I5wtDB
wutb7Tt3FYfOuPWMu+Am5uKBFNiVIg5sVli5ZvYX1lT/L2rqcHhtpSAHPXuHarVdBQ2jXQhNongZ
8iFB1ZPptmlRiGkOXvkxMDbaEcS+ytTirfnsi/jh6JX+3v4ngPcbgd8Lc6DS4X3PDiCOLrHnHN7V
s9RkSwMkpwzwWNzD54/THhcR1eR5XJOG8Xk1NuDsgHLvVpntAwjaEPZbNjMkyFfZc2/eDZT+MQjT
d+tI+PukdbgqcvoktkdIYbNPU8i0bZgnuKC/LwN3GLsUdeodS8iTbZK2MjSQNnHyyTjH5UGOgxjH
rL1b/HebqEwHV3untpo1O9zJSZotHM1dQmzupg+5trmiV3d6UprAHcQ5jDcaEZJdFQeRfqp0aUpN
rY5qaS/VI6ucV7C7/QbiCnRDpab1wfEampvn/IuIwrUy2b0cWiRhoMIJn03XD/P/HkcwhJ2BE3mn
xV87C9/grcg0jnc4Pg197YSml9lwbvQ4YrE55jzv+d0jd1p0P2Z3qI47P1lQ68VZ05Ki/04JDn78
qMgrDZ/621QZFNRhWihmfAYoa5ymyZMG4srwd3fchv0mcUE9cmJj4DKBegPiSXirtTmJGojgcaMd
TDjJ+IwHKjLpKCFFDmrzNij4qYpv3ht7WoIL7/Kcu76/sQaWZLhLB+Uc4LSPQ++/yYePcP3IegwK
OYmPDXuc559yLYvxdgtbx+KjMoLG/OBhv4rCiWGtNA8dwuekAk/L0QskIlM7r9rSNyn56oCCcwM1
UV9A5j0FzORQy8LLAqcrL91ekiIwnbyE+MQ4TlOIfPaevdhWOwjgS3CAHCiCYhLAB/Mv1Nqpb4+G
QKQpIv7tZgdzriopiRIQpsN0rza3nZ5xFbnpyWBGq1BYP3Xn4GXvkJhZZaiYk59L5APmaOzR/1o0
/VfXhKcAPw+JZL/Q6rA1sLct029OeQMED2bqN5fiK/ZjQ7VVYd2ZR6mF+QjZhW/lMWR6XEdd7d1i
knjEMRKZlO+NBgvFH54MlDi0fZ6Fz0wmbpuzqwHON7v3zEGF4Vgo4Hdib7NiG1qsi+RGGtN5PT7L
UQy/wAQGnWXp7aSCuX49u8/ImoVa2Recuflk6DI1BrgBiRWAC9kM1ESBem6xNjRuGCg0t7EoofcK
NLzYQ1ctvICP4n4QNvKEN8yjx8O+Bg7E2cDn6BM/4deftbRQYcJT5lPW+KI6XsT31OIsYYuIYysA
VXN12HubnVlCgRpQzSo4GJjqnwOdY5e4CRsWOfdVExnvSkm5ZvmvGLpI9YVJehdfq0Z1sT9e/mJC
sCJhJA3QJ9FSVAJmFvgLRTACadlr0zQ03/pnYyRSbQaUQPBkRMHpU0q25Oztp6t+eTrdDFGSvVrV
q78TFgMPquLP6fg3gyFQfB7zMQzWBb2R+FxuJVRn/JdXhWjPWq6VNpzB1IAsC/IbQVvZp8We0T5q
MxLqj/EsaHkhoCgIf30jPuZuiK3P0TydvwLmHeq2CnBhvvmVcctp8aDMIhUUDgukSnIpr/VsJI1f
Dd/4BHeRHo/KgFYh70+aNYgfDX+0diN2ofngaBzKHRKGNiSv+hpS9tIC8EOJfVfaRq6FiD8kLEvO
+8vclyZSckWZi9ACCrX/7MeGl9MS+TxAYAzyRx8Cc014zYny3JzgX01fJGGUSqeApcxuDz4Bvmxd
TpGXh+zDMEJBynid0/tlwJGhEnmI8qKrJOy4Og1iX8clTo2stYB6bTcDcDlHSf06+XmKc8l1XuO0
Ljn4z2bRyoZSmLSmHZ3gcAOMbY6FlWdlwe1/jr0ZF5hruIMG3Qr1eS/tCMshfpfIE/a+8qPoHYKW
3QA9xbdcZyFPUpW8CbHNFnHdGlyvLdcJzpoHB9OwnDaUyAMrW7FrzixiBaAr4FfDryWf4nZrPC3d
rueuhohpJYtlNAc0I1P9XJQ8mgXkMosm6DtXb1wjIXc4vWdgatlFTDroSHyKsoiUnDD4rvO0FZL6
Ehni8kfvsfF2pew+zSEtCDobLNVFS3oiHUSm2DjEYNuvETizUOgz0tEvomNsI904CLqWB+drgWhK
T5QFCT8xUEqnKHHU05gYircYV13908yw/h8xLTBgixKd1LKDBt6FK7N20LAi9Ck5BSaYAS0ayXkJ
Q51laElccBVxaKnv3rjC7G9qsrwl+gs62H+/fd0hC6eP8Q1eWYH7rzsRhzzXwZsZ/106Jn9Jf2S4
U1IudvfNez+Pu89Ii4tUSRuVxehpwwJsR/j2qEL5wT4dNx9oZ9vqDN6IKCfJiydNXbw0UfnXhr3v
T7jBPrKinG7Xufvdj7LfW3QhXwv3gv5wZzJO9uzA8XNUt6UEcdHcQuHB5Tlk/9LIP7uu/UD/G2gj
CmLk2TZm3h57kFuPgJBcDr8TSMhVojhHsVtF61M2g8TQ8k+K/3mhGwZeUQeQwwEhJZE4n0UJmEP4
GSlKnSa04+RwFkrXw8GxRX7Fk2/omxTxtnp3wsbVXg9R9dCkUcVS5TfDkLqLTASFQSsDCkEC7z6j
Y11rrGDlPCb7qBpm0kLVZaGv6rlsvGPBx5iAFfgzr77nvtBYEcIGX5ThJhSHuO1gAVCBYQ0+195J
9zMVFwZOGkImgnUJqAdeuUnf5AbAf7pqOsCK2NUc3mINYJCA98Lfb08hrR6LEL5EP//UsXLhU+mU
kCE8U5d243qrm8iV4wSmUrGGD56weO8HDoeSt0cctWwYWKKmPhrlUEzJHZpR+tZ3fCG1+/Ny9yhT
VvUqUXDI4XoAXX38ZMDnFfVKxLnR0mScq5erBHLtOHWGDEcmkP09cJzZYC/AyP2j9on4okolzCNa
rtDxrDS0QH2ALsn0JmclbvqOSy3MqjOZrp5S5A1QlveYdwHrcmNOfRICEm9LwemsAjsHqbk1hYSl
fxZHFrfwg+SkUwM+mfcZ/MR2gQEkHDKz/s3oKfnd46P39abseZ5hr9JzudMtCCS8U/sCIFh9dWXW
WjGVx3u/wtGavqbC5KGsxTmSpVF9nDMVo6bmElhJUBhYyoMg4gPOZeP3Xe827jZTsE0mitiLrTW+
0okfeBBrbC5tR5xGHUflBx0FXjB/1dMYTA7MhFrLV8V+0CWQ9oq5KooLRzmEs5REmvRQXg3s5Gxj
B7pcwTUXhuv5C7YpIBW4oF6WKvXQO3iW+V8on9bHcN2fUucUsdnJl018cAVgXwo/AHylQFk3tRXA
/YroQHGBqLPXEGfW/rf1Qy6YL+8UOZl6x+Y5xYDSYqM4r9rAv5EsCgBjLDWmlWvdLWRT+x+/4ZcK
ovRNVREyAlEkwJFM7NWYxROcjkPcQ2511XFI0K6asYpuY0sZGle66mieh/Lk6a8OpC5oM/nlUQXY
6qI0YAszmpTIkA6PpGvtPN+W4Y5cohtVBjx7byvh8tgBNYcLEbePDLNbkEOA+OKpDA7OVfIeDfeQ
mG6P1oxzYtDOlMo9aWvKrYGs8taYALUxxlAdx6efMXKUDoxmUgY8LrWVetX9lzNRy1I862bX9epO
jrCDLEUTxI1lQENeh43nzDfMM+JqNG5Q6o7bksN1Sa0/4eY34wSI/V9GteVT/faSIow9wuMoUFtE
+a/K5iMY3BmvOsfr5rITMOOg9F+bmvl4QBpP8u0dYNtYDWSrv8UIXFjI00TxCuI4IIRBtU51pnAs
RsjP0CVKTegVMhu8UpuuS2YwD54bmYtzEdoqDC1n3RI8+JbRBgFoZAcQ3ySFmnp1MoVXhu4awMOr
n8a+Ajj0kzByVGNSxM6MjtS89ICbv/e7Ivu+7EHLX4k4Hy6HsIJWoKpO6vlmfmP0++fZT3baYhFU
2CCmhvki5y90FclRQt9evVofyeotbqIFA/CNmOp9wes890JnVrXu9SBO/fgC7A6O94yAScToofau
fWea5h1cNfJKoZMhsL/i3Ln6QIaPrO4pb/nYc8NgShhB2TJX0gvBAqbx75iPYLDGupgN6vn4QJq6
/Sq3Lbegs9baNNJMV8eDltJPj7u+rOsaSPuupHl8qP2cCzq3lbU1oHYZhx4HOrMwqZmgll3pmELg
KNravlurpEn97jLpmfh+jubVpl0DmVbibLiAz2LZboboc+cXfT3nuB3NiQFqIGzn0bZd5sx+/IKu
QuwxGtZsbZjdzu8rnFwQYCvfXqIU9eShq+x/SN0oHuBSUoNYy9u/YrtNfbN0uBbUKQRWxJhqMHsy
OjbHpEncrsoNQokhnKLgZ2wR+HGMrDMdVs/7a7fSO1+K4b21LynYIt0UZU+G2W9chidU1hztukuv
XjbjfKpgA4KsBQBIx91tCr2juSt9OlaG1Hsn7hvYBMe3x61U66DMCLufW/w51BlTGA1swviI5Li0
Re2heIx6tPyud36X/ae8CfC9O48pthEr1ABL2B1FzjY1I9RzULFmfrV73xRYsM4YquzcSTXVxTaP
PF9jDzlFhJwsELkH+yQ4k3XdEJBCrQvEbz5qgb8nGxOh8LQFgoalhCWEtU9nn+kf6Sf0c8Z7hPRr
VGwb7VjALM6lmYOsAC9yO1r6HO09MIr5zTEevMyQA/ctTmuL/nMx6LtMvf40FLNc/DMuTX77I18u
5t1ktfh+Ne4DqbXN8rk28I5pLECgY7vTmGi7W+5GpBt3+eUV1qZ9rRNS9bCDx+KVAXiuNMWJKRnU
oioJrrtScNHgOBw2Kf5MFt6241ca40w4M/LLBr0zp5Tpb/kH8y6GYh+CpfdcvwR7MLHA4yAxCVmM
FjA4xXDjwQNdi7bHVqojwnG9IUhrS+Di2g1Ud9dEASySXHe3LoGiDNazFLp8bq4qcBNirLjP4G4l
C8Dr2Fi6QphMi1DkW0mrkzUPW5z5UV6NkWURJaaueDVA8rqmyWTcE815kOnWKsmdjj281HCugpqm
aHcHzUSC9FLnYyWdSRwO1DhfmVWQ6A73rgxcS8V6tDvA+7pTiPS63M4j6Vkxv3ua3HTlQM0fSTwM
Ga38dWCuLbq5vkeMiH4YhieYub5JrDtzegsSMkP3NfyJ0E8K5ZBe6n49E9XWd1po9z151GTM5wpx
ERnH0MO48JC3dwt+ULQNHSAgqdBbQ6I/fizhrfStW5Sl3dWGLiOu/r7nLpwQj8JXU7VC+O+8m7C5
NF5JRuLirnDsJiAqANG40LKYctPq7YL3H41uLl5k9lcCYrYVZBaZvmNEu7w/K7ksrcama1fCVEAD
6OaSCOv2JpIKQyB6gEY8/ga7DNB58oKNwXlKhijr6s4vl+NSTlLiuHW+ZlbK3rJbtXZbWuDCuG7E
1kiHuvxFEyoAwFJrcTvltdS4Vq1ZwqZesBqZ4bKfsBNW3OatakZSbNWAd60HxjxlAZ/HzFX4TaUU
PNoHZjCAjqEU1AQAY+LUVUyjG7S/+19tN7eYVgZ+gS9pogWd+BvSCGBFrq0vmcZSOTR7dQnFVVC+
R7czh3NmvWW+sMzaTCVNVIELIiCUIY/weBnE+arXF8u7I/0aRfwYRgBfEcgVYfnrdktOeQmq890r
6pvH7nkN6W/jKPJgDFUvjPYdv7pxTV5iNQ4nF9E83uES7pWxEXhuJ8nEFjuVNiaNLhlmkiUEszLN
EYZjn5hV/IavqsTgTu0liYShZvHsbIixb9z8xPOIPGLkdbDxR4Y+sh8XtsxkA6OKry9EXfrl1Ewv
wlBH9oT7wwNO01EAgGrU+ziVsDESrxbSrc+BRN4cFEsTBPezyxLgxEzFLdAm2+0vvixRe95AtSVh
gH7NS7YjJMrzhFz8KgRFNuHf5JOb0J2p6GycRJbL6VbIvDHtpBkR7oxcNTtNwxdMO4EuBtHITjZx
cjLK7E3aWtAcmH5IH4zAWyrPa0vCmrll1J/CTBHbpRYqrdSZ8u9sxYlQWRwdGuz+qCyHVCjN6YDL
/MrCT5lLxbtdnLAaUwITUclvhv06YiAFBWkhZ3bwNMap5jCBF0t1XBMAbna5Nzda8hRsodIsXtfB
0UCOONJ8I53UFN549KEVaPgFpXSqaALpj3QyMdexcSb3/hGAbfWdvP9sNDGoSi4Iz4UgQgHTcOdO
M3bJI208sQlq4EhMg1D1MIWfdqh2R/u8dsx5yBuCOg9mzi9b7HnUz9Bx5GdY8/RrTk1ZDnqv1Yax
1+9VGPiCYaADOzuKCYos77vrD0ZOJukRbxb8o9twGGSo+Rm/iporHFzDxFY0uDaXbzQXEwl1aVaA
hOhs38fC0BYViOTeS+eI6PTp0gjqEIWw8DaD5Pj6OmS+lJexVgm0yqp7yCsvN5ZWSbl0RZHnkqI9
ir2ucE2xbKFozIjgq+Agi+EWvvdj4OendFnVgTjG3x3N+6R3m8pPw91P3m8J6fgfWKM+StYM6Jlk
cbEz/o9ufgPkkxcBXYz5Jg46CzDvQZuexmjioLPwulHHFMCdX1arirBhHmkvWg/C5J72CO1w6KK6
v4xzuZVhTUnPomRuhPR4l57stYoceiVmeVglnDST8ZBwdbX1b3/RD/A8r4PCxjgNzbDaEf+kGzMg
RgXt090EOc+R7g4xPj0+/yZNUzzw2o3djAV86xPgaFYUZzFsFvTQlVfqI8HFOeyfmfBtdJOUwvCW
n1Hhc9ieX2Ceg+q2GUIM8Te6zLqJ32z4+CDDk/W2VuAyf/N7HaKUjY/0Wh1UkbPEu8hHzZB1r3Oe
uISx6t4q5t9P4xM3d7z8WZQyiy/eO7T6DbMxv//HwkP+5mf6kZkYXI/fj7WZNKn3Waij/R9fHy1Z
tDAqlosr29MxQc/w4AYqgzmFAdoAZpf/yHCKYWip8Arym75go5nhWroRW7Poc7AMDnGfTVDxUYhR
OYU+7dB6Di1X4WaWJui7hUjBXMeUA5cVEoweO7ygBj5ELDHHhNJPaRX3ldB6wtL1a0y1DCMIhQha
lAX5dpdhz/LkJ+8vbbF6uAIR1cUs+EEkK9CY9Al587HRpCU4btneFxdR5Uv7/A3FD3IBcMmMy2S8
plZKBN2cz+AugJcDKHf6EUVHZNO5vV76/ZuKHoZeTbX4HsM5c/Qlo4FkaiJ11/VEVAwloeEAqIlj
HyRwTLE8O00g8+HRfY9ATc/2eJpasr/O8/8Ij6XdiXZkogF+G2C1hI2D3Q9ctz0k1zgGGpoHqXkJ
I+2Nazngj2i5xIFSMDF25gCWtQD/VNxtMlPJqwOQmUIVqnhREV86bv9mgYKxyz1neLams3Om0Ip3
bZAJqw+FDhrNNuVMX4JtbEDoGgcfxpuYxKJSaUtYTODiSgmxRdUMhRWjd/F7Ce5mxgJ3ez9NrFSi
cXF/kcUV+pUHpqgYys7YPwS4Se3Pm6m1VZbcwKlyTaAR49oma2qknZ5OHqCL3yCuw8yYt4NQxX+m
G9V28j1THTxflQMNagrF2qpa4pzbtAw0aOiVYn600s1eTWempz1CrAAmEB8OdjFMB7QVAf5A275m
M2wRdZ3HTi0bAF8Y1aE/I77IYoeluZBiH/uu+/X1HsVleX17nGltIeagKKx5rUxTXReSqoRoeynP
Fal7s/LoLB21zAd6ayhtfHRdKZbkVUN+2qLEzVChIh8PXrAZSn1Ys5w4NqNhmRN7h9RgP6qnwgYq
Fg9+UJHczyKRT1+SiBEaKe+xxhJ+PQHUW8HfW4AN+EStSv6Wa/Kn+SjRtUl8rTD2dDRVJiiZfW08
991JJuMZvZiVG7CiaU68CZkxPOyJg6wbDKQ/aRbXv/Am6WXsW7dNFCnxp8YHJoIydZxEawQiavp8
+wD/psKucb92iH2SW94Rb7XzdEEPSNal6NrSDMG9JlWrG/6dosTfc/FjV4y25ANgOup4szbvftgj
z1Z0QFH9DlNQmBNjxLJZcpRHHyzciDy6fsVZJvufHvr4tnzCbcOEFxP7Xjhgu3VB2cW/P15SAN4b
9Ks9qCK4Tq6zCOVQQR3E20lefIFQy37e2vXwgQ5+cMxROsFLykZfEu78KCZ4z2rs1NDxImWORjat
33tdZRvgnJa+Tq38hNvowrde2FJ0rFy0OphvIFID4BXv9BMKEezyUs5QiEKQf283prCSEggVt+3y
bGyVB2ZzYP2openJb7SUo4fbCvYcNT2s6Ato3HAdQ5D9fOkBh2J/KaNFTbKuUi8a1TGEqWuNbJCp
QiGq63RMxsc0IIWkz+Dv/5N7i3pb0tJxSwWwCHQbFG0VsfPLVlgzfC2Whxu0nIxEjbi0Tx4yx2V0
S+jKnia/+i8VzBsvDq1GXHyi0SqnItPBUkpvCeiXnPbw1B1RTsImzs0iB1LEFSj8Oi5pcEbyBmQL
xzr03liz4iFPdFtDA/0PtBFaYrZ8ocuCXsSpsKhwVogKfX+X63JNbavqJq12dL/KZsIpdspngxY6
q7Ce+Ss3FAsSL7fTAAVs8aiHs3Q0hqYogNDXk8iYUZzwMStxQbFM4JAoPlJejcX+1hoi+a79mj90
biQJHnJsADTib0LwXdtsxsp2ZDvhhd7tC5EsuMhnS26yl+vVgB5x8Ycue8Ht0sKomZWh4WjBmWmr
AdyII3CDl8X/KP2ZGrR2EkKgwGAQGnFVttV1elIXa0sgzZom1lg790LlQznNiGacfPcfsGvoEXsi
2AwHTKQp4nHWHm78C9llKapdY06jWUXDwGbYsYq9z/AqEicvVosJH4NqY9F5tOwIoG5H8miwcQEx
KdfFG+mu81ZN043yV8xCLVAP0FYYZdw32OlidLJvyY0A/xYrONc5ux4o37P4n1Wz6ho9ekxkIyuz
rDoxa2vsCXozM1A8+75TP1zo49KBImu0sFUfzQal4ee19xAtFKzU/bfmz6gE3ojQW3DdO63+jKc5
0PDsKC1JRiq5Siq5u7e7rs9XGoDQ+hBxPMPADkNWYsHk4M8gnP0iyT32BCcW6NcOIKy0yXManCl5
7GiI8C9Oj4cpEnrg02S9KekZRbNcmogFaboydAKI2Zi9cJj2DRaiixfeXZcYUojQKk68fIMLA/36
JwzbJ2st1Vefw+Qq+4BTieuBpM1WfAoG5MWM9MCeuEx8gzw0JyhumQhO7IT0nF/LQbOj52HlPT0z
ZWqLNRxJO3BD2aRmoJrt0hKJMIiKyjlVYBB3UtRek3OM1fPmeiXNBElxWf1oXx+4cvj4tro3O67M
MfxM7g/nmbLgRkHADPSefnI8/NFRJDtBgtIy3u3Enb3Bi5SAUtD2iFm0KZv2pvJoPhGxE8S7psIT
togl2p2D5nXNHPQwkxsHjLJ9PXiT8OVM2/iXPwHL+25LeVRNIuvKp8y3q9DlrF1t6bT4NCUYGHd0
9jBhDY/0RiRtxGzeJhEhki9ZzPCCffta++RIytj3u9erf7iUUcFOUdyWOg2K3MvQXCw9t8dL82Xy
3qig7PbVUtEfyyMJ2jXVr9RlPOlV6CIa/jK4YcaOprl1W7pklcpQowq4jL4M+//CkZ2TyoOHOqJu
P5/Wg5uFFJsRZa/pujArkcbW7/rqeGqHQwhFnCI05WwMXN6XLV7zXlG8jz/hk/ZZfG2ghR29sySi
JhABSTiMZZwGcH/lWF9qLJXMCB1Iq2c5abZ8JRUhI21bquKJbHmgJWzPKq0FLmWu/yq21TYDIwFG
F5UGc5pqdDR1g4LqEBGk3KmBZ2X3ubAJVf3trJy85SU5wTdAEzuQeTcqiEp4gqP9BiSfJ6ydhFlP
mTpx5DyPlJxnscuOfEYrjW1+E0kWzSJgSnp/AWIHyP/DlC3RC0B4Et5oHoMDjeX0o0hHZd7pAVkQ
C3o5Qk6WOXS+RHZtK0ecCqVjrW0LaK3TQ2B6YWVH3U8bz4QLJwMkC4bp/bHun2GkVI43fE3LgP1S
S7doVcaxUAcshMS1uinlB9Lxmksfm7P0U8X4RHM/i7mBFPAQe2RRAxe5H1dIGx1ca9QkC7BFHbEB
kflXFFPWIvP5HTiT49WyuIdbP6VNGyR3jNI3do9SqkapW9SbZMfb5CpeWIxxA9reAUYpodv1IT9S
Vpq43b28OUWGzhOme/k68D91i9KJ/H5KLfv2n82vWnv2uD3tLsrcVDZ3k3vWeHBLf836jTkwNeGs
+qaTcCYjopCjd8UcDcXkeZi6ruBs/QioJaP8RcX9jPRByxLycjYSeWELJ0NywteA/i5+1mP35NOR
CBdgFYQv25NW5AtnxSr8OB5dFjjwKThJTVaOO5dfzMuhx4ol0GrpbCKI7Ml+zPkfx0Ser6TGIUgt
B6ktieIvGvw7oKfFbPD/X1wl2ZLYusR1hcH31xVI/f2JDlc+XLbfsnr97xBWosc3LX3Lx1IeZrtf
sTs3ec0U9neyGXsf6jeL7no6S1awA4T9kfYmYlDQEUd0XJH58dLkdMa9qK4S0DznONSM6b6pT+89
Efq0oaGmVWIifWJWcTr0Jm/cr9/TCKbLl53RS/txQ0J7p8KVLnu1cZ8gDqZabN4ypOMGohtxPiPx
fyJgjHHlfBVYXwjfZDEueFmMdxEWI4rbPy5aSGxYo0jbKP9jOWaRgDYon7JdltgjQ/fmyhH7B5P0
KKcb+L+f4zBxnYoALEb4IX6Z1Me4Wds1UYEmSTzB7NdZwZ3MGO2140BIAlw4BAGTjo5+ZpGcb5ZH
0nzLwgEgOmWIcsqu/cKeLeOX20/yBIS4hjvZrVD+JTNE8IO3QpujEbMX24v7wETCKFj6Ios0ZWiq
FewgIIgYbO6DaWu7Ts4xVEN7DDk6dOG9iI69PrALKCzJCxg6bmoWOzd+jzIDvx0ULFtq72hsqYix
Mhzz1WjbgZ7MW0Pnv46zGxAxV1BhNuSjiPuUNHXwRPTIvqo6KTuHmCKGnxQYyPtd3wOvn8hWzKKU
DNJM7bBm17yoEXH5AGM6mYtW+mjUTav1kpkgpVnWbK2RsD6FQwKLN5gBR3ncewEgjM9FcHeENXqU
Bd+Ody4omkIBhRZbX5wuaKnnUBjrDvj/fstP0/WzTcemKnsuySwv+QRqZAL2ubq4GqL8TfmrsVWE
RKd1KgR22UfagkA/MSWqIMv5oRPsiFBwd0dXHc37f/G8NDQr42VH1h7qmMT2thl7wpL4C8k44wID
mPd7Yli+k8uZJjCEL54dK+4TDGEMs8BOGZHjmD3bX7mBYB42AlORedWed4zNRnu/77sFnUFb4Yk9
1DviMnV3Mg39Y83I5Rik4Jj7uXS1z3LruIH7veq3noyOiYXp1Xap1WA6EukPyBSdhy+5iMZoQdaT
bHsERAwiYCdxVlM3LlETCt9fVUDMusMJx9BLdYqjJzkGysTAQ2BiujqY0PjxdJiGnKJercodSOom
7Y/ZdFrxf6BBaAquAZsJjCAp6eLv2DBdM5cG5BLb8tl7r/CGO1qNSPcaVuoLeAlBuX74hDfjQjHo
iT7SA3pLTlwFp01UOTZQiEmoV57q+ca+Tgjj59RG8pqU2TOmq6eqT49Cft//uqqHdvns0plJGbp/
1q0nc2O8flyZABiBvJfSMH0RR38Wijy4UxaAUcxnzdsFFE6pUg+LRBMQyOJ0pDRJrPWVyF6xxTjh
hSyZfjkm/IJyMfz9bKa5MYIYqwJqA0+gRsMUbyRqfbVtF+ZkDlkQVNf1cRWNagd3/IxftXht2C5c
QJBKvKwy6gxj/g8SC3HV4nK6vHF9nmJixyC1q3wSJWVdamSipAPZUxyt/LyP0b8omY/3h1w7+24j
Amyi3nNU8xL7bsSzb3SDW/lzV7SjMfCb5N5ZWeA3KZqSLs3s7rRuhSxtXL+v1eY7lfdMbA3vb63U
AQyEfOmIeV3VLhmvUmA2BYIeNJx9mybzkODhaUwxLuhWm0NsMRITg1gWp8tI85qePJzUOgwow/g7
AhMuBcSNcjdz/qj69bRwA1gsfK5QIQwmojtE4aFJhZe/YBQbPIVSk7y4azDPBA+XodqVnp3qjDaR
E8FWd8/FB8XuasvDUR7EeOiLDU3URAL43CplcKY8fs9tekddyBTF4GKrncKw9zAXLR9aH0KYuFvE
OkjZjKrZTgLngsfngF4+TUNUf5RFj6t2eL80NUvyluqvHAtMX/Zhow4gjVfjf+oOfi2kr/G3+uw8
5yR5Q2fcdaWMOrDJQNlGbdx87NFvCbvfQOvntug7BSRVqHfr4cpU5mgbsiEdeY6T3vBmvS2HymLc
in6AeFiT543w67abPaASD0ai644TE6i2tA8rq2X5M7udu85Y2a2ZvWhnX4Qh/kpShAjGy0CPLjDt
s5wJnmH3uBAtdrGnFw3CMvMKEEqdW1Rrr+1Kig3iGrSilG78+ljvh/c+Jf7TyxrI8S5lYzzrjo61
FBtm9U9lFrypkHKfQdMQnj/8RtvFhBbo+emXA3U+nFBarAVCzds9ic86oA7AM5EvgBuVvKTBC/cq
1aa4AWlKKKhUZi1TPxbHNF3HqzroBWSPm8Sq0cp8z5xzm2s8Zkna64A1rkT5Bt7lU8sVGIpaJIL2
CuKVH59rCsDIfaNuScJqftZAjMl8rKxxrR64NqrsF4G+gfvN3bi7c98APtQGzeuD7lJPED1Kustp
BktWjRl13aMDdACCTl55yw9kba4HfFpiSqpyfYyVD5rnlpryCTWZaWbIp1DthNLDfUUXXo6mHi/a
oFdDZLC5LKe2tlNsjtqnsgr2EVZ4zFMhdyykyGtXFLyoGIMmqn2Iha2Bwgx7RYKrk00YgBavzU4x
NHebwtpF9JmufUoqSSP9Tt5wNxxz5vAZY+xZ+v7n6vNGzm4S7+Mi2o8GPjXp3bvfqmKTuZVcEpSa
+EQMSxRe6ydtluz6oCayiEHfXKso9/sxeiJ8jBEZQUPc8SYYFav/2xmTXzIJGmc596GRFdwRiUu/
BXa/RwRbV7FwqvEulC1CqSJub/iZGnjMqCeECpojlRdIFpYCDLRuJFs5SbC22ETS4PACiv1yg/1Y
FfPNalwco12FQwg1M/yi+rEpKLxLxZtbaYwt7zfJWY1Sw1sIH00JD91eID5S1VHpnoVuv1XdCG49
6K0RSkivmg3IeTCJrmq0llCfwYP1PlXENTIMLe/CaPjP
`protect end_protected
