-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
RgpoBtGJ8wvbTVQop6rnqPT1m+RM4Ixycnh2mssw95EUxsgb0e3sc0FMRJRY8v+fqKREnSzIViRf
xUcih3abCsTuk19p1Sx85cfqviy8Kn9kFflBIZqdp+4vNRpH+AWAaOZNMuj0H1Q57rynipFgkVfz
LX82P0aH7nzxjYfI9mY+Ax2oFFwM6WJB4kXptrUkXd/fN/crQ3u1LDWSfp2V+cGPdZHx8qLoyRCX
s4MsDnsaI049WWrZlAMFdJ3Ghqj975zb0UBzCLFdTKMi4w8xscJ6fmNYcUsmiMxC0ERGVDgCwuIP
Xy9I/pBcOh0PYSld6YgX4znPxdls1bcFx5FU4A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 24704)
`protect data_block
xcQrI4chwP/GByYQ1cbVNCbiDRp/INk4fAOS3+0NdZSbLUHPx6kfXpL+Wwner0JgtGq/v+VFHVNl
cclM3rkQUD9hL0ecmh9ylfSEX90jzxtH2MkQtqLTXR8N7E+g3Vi3Yu6oYDZZwSXYWP1WhmL+MKYY
WzlPlpc8UY5onokHFwNNsCixhAZJFsGlQPMNW9+Ojs2mgC4J47PTE7s1Puif3hbvI3dj/pQy2ybe
NYFVPfKslk/SAqJ8G/9DQGH9l7te57/ZU5e/zuIprUsOdPeb7V/IZLgb0EdjTFZ1baVDahtpJcr6
r+K4MflBfqv4q9mlsvHnmo8QoS+PVducgoYL4izbAsjN92ef3aq449eNXMQ74EWVVFyT/APH7qgz
Cei42eG2Q6Ko3jTz/TxPr+FbEzXUfJlXn6eElnPfbNWH2pTDRSGPiZ05K9/5wH1l4LpfEtPIEm87
UnKJolpQwQHJCrOTuVqaPgv4xJolYI0qBb8RHmY7z8/Hs7q8V5HcDQtSN8vRRCS0WlzQyaS8LHAq
nKVWVSLM52t0K5zRvl6Xhxi7IrvT+GIbKduxyHzaCQzs/CWIrdqOafCIoetvJmWNBd/HJUiXQ0mu
5xjizdtvwfDr/+XA5trBnzkBW1j6A7MYFtajouJwK0w9KCLc0Vz7F8wkyEV+GeL5dBiroio+CyTL
cj4rI2lNsuW7kApekru1IGEbWrjsgD7lg/BSj3HJXfOq4YLaGkly0zXeikloiGug7WrqYHEKlbwT
H3Exdg8PTK1Ux7NOqld6mW68rmOmKEGO9uOs02Z2AdFTevwaaL0tpCdii8uvqYff5hKSKNA20sJJ
yhvNLeA+PVCzJSjGGUybo2DgLfyvviUdta2/jMGJoxJyT5eHZOsMmCjyGVjBmveOqIOD5lRe0R+N
k7PbNUtRGrgRBI9s/yhEVKkkYlLqeSy6L8KMRE80TW3OOfDWklqmY0MGPbMtB+0KF7FKxxU2aVl0
n4k+Xp37GC6H1jlZbdSZ4PjqOr2YfcfvVHr007nlAKtbUNtaf6bLZfJyILTHOy2+DJk0M/TNbY1q
KnIr9r2tteATiOa0LLm1siSVLrayQoMYfG5geN3092RHw048oIMJIWT/TxWiuk2iF7FA6EC7WehA
K+lIgpfeicr2yXG90j6IdZH5VQdCAiW8vYRKdHl6tXgGtEtNelP7DxqUuNLdLdymUFy/E69r9eD1
rCC0ab8eskaRRoQbwEXYiwqotSvO/M7X5Bl1LZ53MbBc1HHf09OwftFX55OhchzrrILokiivmx1Q
u00upDd2TqEZ4+UyXPclxT93m9emvcJP0b9mfpMpPAjYQyOlWYczYOV5Qu7RixvYaMtuXe1YSpxd
4Yb6Z4dAl4IcLNdCjcapO9vr61Iv7yk2a7HcasHwkftpE4Fdc1Snf2wgCKEgWPYRgoc9sLl0PaDl
RU4H4gl8kmEIQdUN4kQxsOgtlqHTSmYckw/NYdIQY5MuwSXm+9d23eNtNRv2ONulgxAJGzq8VV7Z
GeEj07NGEzV2J80gY+GVIPJYKSSuFh93rSUQ+Eiky/LhbMLdFxyR9Yeuufl+19VeoYNLzp4BcBiH
ah/HSl0D1UUQnzA4OTlap7mQuD1LuXvtXHMmpU/HMZO9rSUht/DRhWGQzDBjHFVPtaWFj1a4CHHh
Zwkul3AH+Mmlk/lv5hK3mVxT2zrb7pzYLklbuLP3vtHY1cUtpk0a9Q+X/5/zh5HPFjWH/Uw2Xwjl
Ss3x2+lZb0myaaJysRZPn22SRemEOpI949loSsNT5ZyfGLQTVnr9hWFwm6m7KwPI/tI7/+gLHhIV
Uiw0LBMAF2RX+oMOiSCc1joqPXyXytETpGCVJ7PYONM/OCHVLzmfj9+eej9pJfYDezmiSBbcRhW1
6zY/DH8WEIGpJycPptprg8U/dtBawwYNgcqKAI0ZWF/6za6GT9NW2AoHI2XyzRDH6HajuhON8NzO
ktT1QHJ6/AI8vVwadxVUlzTsPpgiRrKl/o26QKDgLuOx3jmFfQtFbJLD75GB9ymJPLXBvxN5iAq0
Xau2CvjlvM2RwnemfIBilnVSqAB/UWM7fpLaScM3Dk6N/NKHZnNL5ooCj2UISaYaudLoGv/hewuq
ID6g5Cn6bPU4jALSMGJa+EMv7AUyKPT1zscn9j0Nct0v2/0JwBAuOq0YxpbaPvHdF2n7Sa88kRze
qPoMLZEtttD/Wa10PsnZ/kY8Xoda304VZfk2vVXn/644ohq1eRBUo01sZtjFI9+RkcISsSJDMPOm
jlG+VZ8P7SmE0RE9MOjRSnRADojnGJTakY1cD4nvd9n439YhOmYSU18q4LTpf6evNDAM4MlDhIDX
dMoHLzO2ax7GPX8m55HAfL3VPwxgVlXfgGTC39rsYaTFDL8vajQQjNsIhJCoH9FhQuRg6MeGhDAy
LsAb+Y4D59X5kIvwCttlIAVk22PePvjSQjrXOXtU5Rgaayvsqx1mufBzXgkCARpn57BxzIp8Cs2M
SM8mZQuSayEbABhpUyhlhO44rs7ElLlb8cMfbbceY4iiZMIQ0gn+3DG9VTdryEkpF5Au3Y1WNkBU
Iyx/9D48IJCIQmdN2rcdHgfKRIbLXa1p354FmP2S0gBCia81+6AyWFVFggCktdiu/okWc2xeFOjK
mwS+gk4+IXY7UvzBJKzk5mrJNAQP+Im40OM+oGESAlR1Qa3xQrbni0PfujHeI4Y+D3L5roVhHkQS
qsQHqNj0ldfZmGeaFdhMCXQkuMxRSh6KZxiAIQlVEh6x0ikjKpeYXsGPBDyAnFmWTcjN20f7uUd0
oov3ZY+TmJUSirOY3WInNQdVbH0iyh9zDCZ5unW1gT7iU0phbGVomEu2Pryeq8rDb/Kw3Hf7dBB/
M9PZZIt0Iartxpc1p/w7vAEOHCQk2kLXRGvu0cOvxEgqS5WLfT0Ug7AgU4Ib+c9JK9clCTLkqyaj
DbmaKat2mbwKnQej0sgRZm7JpJm3LMOEahzpSigXcwXD3ptdakfVY15r+uCJ6xgRaj/NfKG3/51e
ziM2wFplKxQhlKHFq3BUgevtoDQ9iFYsCuxjNtcwQNq84HkCb0GL6ndTTE0zi2ib7mOpVM2oyv/k
jqGIflI7a3noA6NUBvOG4vVHfmFBGm9vX+sGmDv0l0UAT046r33vmpVRDM7ywJJ/B0JrEdxrzp/V
cGT80nCssfZJhJPemfPxMX+4sy3XOOzAzQBBU5ZrxbY+0aylQeLwJ7sEI2Du4slxctzKR1N9tdwV
Mb8S0OHeLqRoHET5TyAROfH3VPa8QDPRKxZU9opkiagnaCT3NVfMTugFejEocD2c6u1y/Mgtyl8r
FPdwlx24jTOa4NkRGLJXOdswxrZvH36IV0/RUfAngNEl8D+xkRCLP1A3WH5vVD1RMtsQeRxtL3Vw
Q6k2+/23UNOK4fw4SsNuxJApmZMn1Ks5PB8U2tFlvcb+LC7NJK2w2mEKPcKjzRnbvFshGfbjrn76
aSioivmTzTel+kRRx8bIJYj4AuckQv3col1kVsGg0h8z9F+sBjdMNAOG6sqrBEYFNJ12iwZ7ev0d
7h2pU231LmkKeW5vI+U1aT/2nyESDUz8aE4aOPARd9RdYVsso4sgX+GFe5G/O5sLlevEs6QNi5kt
2rTpH1tRnRLBhZycfSxUx4J8/KUk0MJBkjJ6+Y25hybWA4TYrYRlUI4Vjy0eaCF3m8eFgeZbLToo
neOqQiIWEd9jDXKMkMzQlbfXLu9i9bsYZX+Wmrl2o+ZQhufYnxMBV6mQLGT2AY9UXY+Ta0xj7v4i
bZN09lExoNJzMwdUoQiwSaKpUI3Rt2u+V2bDcTISizQW4m4Qwxs/4rZ+7oJc3gISSV4emA6DDaf2
8CgtsqHb3YQpeLeQRk63wVFDNF7nS4B8+8PU46QYhcLbIQjkGGnCL3L/2FF40P9ThuhhYNEOaLPk
jfGifGt8RbB1hyYhRe7ZpXH9DtKwIE1Doa8LmJQZiz3XdkcXDPKlNBQEReNDuVJms1XZEcOh0RDm
T4i425C91HgVp9DARX7zA+Mj2fdDSiDY1h/A1tZT5Iqsz5ZB6uQTH1Znh8rmMfVecZlod71j6N54
UURi0tV5gSBOpb26y3c/Z9CHAXbnZK6tjiIsKSSXQND+Al9FYQ8lTfqadD8q2tl5XIFCSecn6XUq
cl0mWVQY9JrK8r4Cxpp0eV0hc2gkO6MZsc/is4bz5PmCMQfYdYGTDxpwJuO4VquXTSArOXxFu6Ti
4iyxEVsBJLoGBamW5WGTtaA8wnKaM/15uEZYjQi8wlLHGOsX5o0cVa/SWP04v2SVhzNyCxyinID8
Dufd6IohjDF9AFvjAjGE2etwkWNme8OEX6Os9oPBIECRc5wNo6nkHblZtjPhm9D+yPV8j+p7niEo
QAQfVE3gBZcv9zFtrk1KEguD4q4YAUfUqxlbjg+n3PGPDX9vQEFdnhtb5kHHJ2uEo662PFqhoSfJ
zvQB3bGuInT6XxsoEN7Qw3tFgmmR8hmqUPpOlbQ9P+gOeKkTfCL6x/NrksGubFiPEHWRFURMwWA2
Anl+zPVKl+j5aY/tVB+7Iet4BTMqKJjnkJdYmgIi7zTmdoS3kP/8SSUYq8ZZDNdq7ZBWy63+OROC
INp5pWRgHr/6vIX0eW5tF4BA57FlPOsYe4D6UNu11HXxtzb7wRa+o4U8E4rzOSL8EXwwKTI0/gZ8
w+Y7x5v7VX6y1uThsWLeSrFnubOexNutaLx5byhW4GvnDU+sPE55OBwxZefcp8xBT4uEpQvuLR86
Xyf9w1kG876ypKsf068y4ngAd2XPJmpz6V9lCFytDHXKnSTOAulXLONtuClZGlmwYsawcnprBr+Q
197aw7hlPeOK+8a4DK1v5Tio7Isdp9xud5wu06wGgSd6D4w3lJSbJuZaSMq3AUvFt1CoC8bPf5qc
dcRYr/GTR/s92K3M05U6R4YjpUuJag5MfPMxBA+mkTuzHQwNrAwWuzgatKbbmQN4Ox+iyvjEkP3i
IpTRSE2KKyOUXhJ7rttqCLvNNIrieiu+AMuU/XPxu42eih2GjMzYIV1BdEV9uRhi40OTryurElNC
/1lOaObNKU5vlVrG4B5rgr3zE0xdkobVb6s34RBLoMaTUlOLlDDk8SIZgbzyK+7ZLj7r9ALNb0uI
kGpoalG9UPWoNNBeiOcVw6a4J8HqyJMHMvEkykqSMIujlOUq4jeXJ7unrIjXPgzoOhZuTGZdcbnE
Ghi8cjZfu/ba+Oq2BZwFO/3S0zI/SCuT3Z53AxH4/XzTUH9bRma7OuaCHbLy9QpdhZSrN1Ppxd1s
w7wIoaQT7PagJeHU26dlWM/qiDOqc57E8g0P8CQxR6e4y4kq0hQqTSvXzcAaG8pJIHnnYpoF2XEB
yFB7pSL5pwUgkkAkRnny4BP4witc/tjb6tRRzuu/mSynIvygIYRzAa4k/KwOogePGDfzOcEIMj4w
uwa5tbLvVZo5kmzADQDNL2gKCnlrr92Q9HIdpyMcO3JYnGngwuwcUEWv95UrrcLvfIb+pa9RzEB9
IfhgufNt5Pnxd8nLGzHHGmrevOGMNMQFS1h7ykZEQfnqlpwtklNRGx+W27Qqmfbb6yiBrfDrHRwR
HSdLB3X/DO71UhlfO3YH8NDRYd6zVH3CPZ+Xa/5OvkUGNGp9f2BMrTUbGTaUPadMNw7a8HrrfTVl
wpXCpIPXbOFLRjh9mnxU8IOaBKH3YznwSTD7q7oPpje6aDgfw+/Jb7ACW62vix7mEwXdWzzdInKj
+y/s7vRNaO2dIJYN+vWRtzJTRXCTk0sz7UxW6TUCiAJ1f0b1H1uPCzwHB+aEAu13PeQR5vvVz28b
8euzrWBu2hTITC8z5MgE+WT4REbPiuGAwAFJ0HolXpP6yT3KlHUzxRBWh5G5VtMptwuems2JDroG
IyuQIk9SdcDKV/FB4MswAK4rkH7JKf6njtwi1iCK7yYVLOVai3ao2Itr9qtqWrVi0VlsDd+YjxRt
y7Dm4pWDDAcX/2k7vbEq/K7UJV6pvJ1j6NGR6qwV09MhGq2fEG3OBnKQHyQbNH+pzVeZiFbTOR4X
V9kBqA3yVtBmoK4PKW9pBKf8iPLfwZ1GEGlrcrNsbRkAmW8jIV77C55blRlvDupYsP2VxM4x1/vj
05pN6E/u0p2RIUCTzoV2sK2xNiX0M5SsV61UCB7PZGQ9IbM2uNJYqZp7woPL4SEeqBBZx8aS73hf
FDFGbZuIp8Iq2iSFzWK1bhfKcnALn1aYc4Lt8hil6seQ/uAz2aK36z7v80GzkyxTnIfy/KUtlqDv
KBsvkFH/Js8BzTuh/8t1hABu7GY2ReWpB7Cvh56DHNIdI0lPUGN/vpYQ2dQwJE/xlkbgV340t+ZM
VEfro1QZUzlqi0EgJFbHAigYtr+a0OdsLZzUK3fG2ez1CMK9kZOjzjXbJc4yS8bh2Wa+ixEVVwA2
bmg2GT4cwyT0U1At1ONhp6dpeHSsH9GWOBP3s565dV8HXLV/7HvjmTc4OijNG92FbL4m4fbQSXmE
0tsfTF2hB5zxIrMjq5XksvA1hYB+0LnQ6DWobgo+QFotoBHNhUxfvh0nuUFEBoyIhDTKLMK7BPHU
ApRAjr42WUcteg9TJyJNhXOf26PntgO4A6tfG8I5lfF0OFan9AH4UIfuVaaSnZu7i8WP39G1gZhZ
Mv9q6x8UVHHdGzglRsFrBzYeRRA2JG4jI5GkW5/cjetfeKyI/Y3PQXTf3NDntjEuVpfvs/l3/GVN
PB1qtz/HzX+lKkuaVzU1+fcDILdfuSvx+N7yp7MVy0LIoCr1WsDUCqKpR2/ggtCni/4DhE2md/ea
CWviZ4sS2he5HzuKJAoTq5xIFjxhAu3jfM9U9aPQh9SU2hNo5AaBS54wNyt/yZB6JyWRSgSB/4ob
pATI+CY/ZP8Og5jmsSNLjbffCcge4T3ttCVjKqXB92fIvHo+T97HAxuEgAxbKsiSNi6TtuyJrv3u
PHG92xr7/0RF0k8eQDt9SZYvSmPlFoSqtwRU8pr8a+sTzxqq5K0v4LfOfhIAE5T5Okf3gOoVyDEO
Wl28vzI+VM8+2TSo3mgBVC8sLybKSsKlrE1OfxrUcH9j9d3kvp23JOWep/tySLxXxx4C080EQcMn
LxFSuyev/sEtRWd00UtqaMrJdOUEdDvJfomIk3HWntI4N6zWMUBZMU1ahQO78V5Y4b3ZR4ujixaG
2cFfX9BU4IVUxt4D2tO6DwnuvQf6AH1k3BjWCYNyjSK1lFjygS4humcOlVbzoxPQMN9QpgWZ0rmZ
2q7v9lG7wIMKOxxI1/4aOxcYRKiuCE9smf5FIBaSz0opIReZq3eTwhWyu8vX6qEit2Y5pvl81cAd
/AAzSs/Rt9cPc+KSrNEjDTW27FV6nqpTHnvWdOzVFSAz5UdeBM+kPkuRB+Hv3ZxIrAlubRk0/rD+
xBKeHwqnvFNhJHFBOcv0T+aeiVdisSAkupWmm75vX0UJ7LEsp88MpO/ZeeeR0gdRrLr+7QFh/pTJ
8ZK9okMsO9gCTmJ9Tm865cDcIkR5l5FRtpYuysdd65vpRMR+iBlJEM3jsOU74/Dftl3Hhaa/AYFz
S9Q9icZta7dkGYICYlwg9tYZ2FCrThX5/OVzIegM05l8aWOUsESwrEA4twAtVqkSwr/GUXIjnlVf
BuwNLVfwDUwkyD/ofsm1gXJkLxRWat8jetfrelz5vA58PHFk/AdTM49b3F8sVC3+oGjRO53ocxQd
ZFa9lTD3Vs5aVmXLLfStJ8bO60+bX6AuTfz55EoP0z0RNMEb4WHipZayzrihgowihmLdAn4MjjlO
LT1+cfV3oMCXBfLxYbyVrXcqScOaDqyfhJBcWcRF914i4W+Z1+wqTRuVkN3XN1wqcf14aYTYOnX2
Xb9Ht/QbXAT7kiP/UFnBf+gmXvfIV2aT9jfqSexMAFM7rmfQzqoA9LSnV/LAR1cT0gYy9uERlaHy
VY6y1Qi93z9WSkzgOKr5iyK5p1nWcRJPmQ0nC0E3jJ88Ut5CjbRPoFsR2z3HTZ0j7PrAD2yzpGLJ
WHkAlpSfFct4N+1HRgs0hOQIBPCIoJlBvvOL4KcCWUnD3NHTNSe1gnC/8sS1kqYywQAy0cOQ7z/G
5W3uNIbIcdpMSZ0mUpy7rkzaeiukr8s2AJXT+B0JlZlk64+ojW5DfZsmKvHVvqxwVkBNhXMu76mr
9gvDPwgsTWdwNQrCe88+LtXa1aCjkizvF+LS4X0WOYfhyLFHOUH3S3BcG3YBrEo3F6KJ4okXGQGI
AAuebxzePWvFt58XLvO2/MiJaqL2Mj7QcXiETKFNEWEMlQwOG3nYBSagkwUv1h2nh1gJn+JrGTwj
HSv8XWnBcTKduCMtSketZGZQEx9JF7IcxK5xppXM6Oz4QxRFf3dx+O5lL8FcWtJ9J7XGQ8L4bbQU
QBflvIf08YJhNXEF3Jpkuk07l0vQEtBaM5piZQy/jCOCM+L6gZNlbC9gW2X2GCxVdIGHoglB7hcw
L+s/BlSAmE7sk/u2xCC5AyHTH7kpRW92mTIUXJ0KggRQXtC8pS7/2ZadtetPmzsMP/OR/Q9svv00
GQdLS+Epz3JZhnSMPLOfOX4iwEhQVQkkmmDp+FJTJc/kBRAOS+OwyJAy/CW73LESanvfNKxUfJ9W
plzwpMFzDaaZPLjWvxk9Z27UDIrk561RyGgy79nCcLELY8tf+By7PTTwA7lFo1vOSEYQSp1lvs6/
h8z1IhUx0ItWwRJnI9hMqjLcIYcYGC8iwWudYt/v1RGTkzqX6IsYpMU8/UbzRvsP+RPG138gzQoN
QNBWjGO0EWS5LxxWhztGb89qJQYcWy7xw6s/sDLkund70ioYQClwy3lCWWU9KwjLEGDlU86pduHW
WB/KzRakQ2Q7oFCaeF4Aw2DXFbANoG6RW3ozarOktHuKCe6tG5pmq4A10+VR6s5sZMlWUXpAuUxq
P7KdkXLhIuIEc8kNv3MVVrrZNVUQX59S5AN9s5a4o7luaq5boP9T3NaCSfiAs8tqguifqiJGgiox
jEiN9oeOFOjzor8u1/5isM18LO7sFe18h1JoaqQmiO/hCsafZq7SSeB2ICzTSs9kZ38622adsRur
Z2fcphsd4sai97Z+6ir5vU3uchNVcIg2oJTsvny55Giq5ClHbPAsp5AwdqsOd0PJzOfYAPsXYRNT
tHi4rsbkaPIYAelAeZTqHCn+x8Oj5lrLoeLriYct2kK1UPMTyieanJZxfZMpOetqU742DXjxe5oy
iW2uZtWNjn28uhYi+EdKLi2U6a4j2/6QLADXep758fTpMUDn6w8r+jENBaj8/cAg72tpFihfeWDL
CyjCXFaMTaPDfRUWu5waZCeUIx2szh23K/ZHF5QLvLqBpbLEvbZVfF7ejeiq8P5UtzYVi4zIzb4P
r014XG+qQ0I0TO0xwDM+ndCJpEukATPKEhzybdWSKWD3jTQeN7fxA6grnuAWkgmKHB2kX4jljM6f
xal4STqPoKdysaAo7dAKViDAN1DIhRUpqyxVAkdvRSZYPph5b2j6f/aWbN2/A5orYoerswdwizU1
ClfGkvkNbC+8ia/UstWZZSzrjT/KLjAgVqWe7N2/3WcS1QWYgNP8wiBRQRPv2qOZvDRgNd/gQX73
V6bt+/jMoXKVNCr7ififA+qSZ2nV4FPtRdMEnE+EhBLLo9qs/a1WlKY6PUldkJ3vLF2QwaBLlLkz
zKLB0sGEQlqDLmTNBXCm8f4ybvUb4HSpBBQWY+cxhcVZWjMocPoz1D+OLnKrGN4zvK9LzqM427ec
vMSN0QwS0O5TLgWrDMQu5p7TKrNvf7XOeMomnU+bxQBWjg0XwdEFSw2oEpW5NuEJybHLedPN4X2o
2wHBn26Uv4QTH27krYEWLr09ZMBVgint3HerkwBs3z6o3qkthBMAgpwsaBh4r1eUp3R+R+bFrthV
JVlTEnUSrDkqm81CEvpuV4L3RxytnFtudFQawDqBvALB8IbiMjEVKIzHT7UAFkp5OHie1BRHimrz
iEBfQSHsQbQ4hJt2PYZM3Hh63UxoenQOqGkO0GnM06jTYjWYpBz0cOrn/9CFlBqEQ20NrDl+hu9i
8LzUT5Ee+Ccuc8r92Wv0O3WeEoG7eUAM3lpy50mgqECwGQacQ4zohG9lvN8EtIc66jH33pUnhLTj
v6sCB7wluD07zSxLcWdmCPEh8kzbDczi92SIs3cl75NHZ0o/cPfxNL6M5xbbk3hnyS0VSIwhu1Ir
u+cylcywm9I4UUVqwk0z73wAYgGem3Fmr0rY5aoG9P10RZTYvy8Et5ghqZAmVHldT5dZcb8474ny
ljckujNOJ1B09UxOp8Hf9R2uGXSc1QcH8NtltXrMIrdylJr0YVyhLTqjwEzmDeggsVgW2ZjbDHtX
8DRUBo1OuB6vOKWpb7JrkhuS761AMGBUi+q3f9G9W5UjwSTEbxxAvkDo/epsZc9d7+DKI+2JB69q
SrSum6QfKIp9K1W7LwF/Qiwy4hQ+uZYpd9pYZpP0ly2dvdR+Did+GyMD9I3QDLmXs+5Sq0rNCZA8
fDMAG2IbeM3B3qDO9XuM1aOO2lO0RYa5iUWBXXt238Lcd/h2H9tAnZrr9vnIk+rV8Gb8+DtDU/qM
gEFxYUDcxRFH2j7/MJRcSU7ds1F4U7Bud3j4fXysx8zvllQ1Nb7RdRGtwMmEgMYovyyvv0T/cfCE
bu2FKaxv/ZPwFZne1ddBGkb+utpKajZtKh6mZ/EaXwfJyyMsUMHe165hCoWgBYmSZ882Buaw5UE0
3Ad6MxvM51JxTC3VUUfVV6dgyE60790mwaMejILoV8J+hn0Ik8FZo+NJh2xsTczkjQurO9/0TLDd
7uVVkENiorghlaLm0WrSoA/2Ik8PT3uLq3CdDoSl6/GeNxn4SrCDqtKWn7LziuDhZl9gUHCU/Yt4
+WJFPPqrbJNgonqNOZVTek1+3FtsQeBjz7jF4Iwwz8YkyWgvQ1sWMR5f2AhWVVQf6TCZ/gsPi5oo
ZjkTtmESFWf7wocMP/QsdZFDU0JWdrIJjupI9Sujd1YprukQK99WRbiLkws8ChmI//hoZyoTrDq7
Nrvxv2kAf4kk3e1zzv8thD02FoYWDdOfCStm2xsIXXHIIh17h6IyyOFaV7SaJzvrSTDNBAofGE8s
N6xbVTlNydSxX8hYXpE5T03wgHTRVj0gnxYI53X+aKq2N4Y5/qrPJLG2t4UhWvbRwjVhA62A9PHA
vm279/IsPmR27nN4R2IGJVQc/UFGU66KZC7JrQ5Vf3n/kK4Aes5kl7R5D10WA1BmIx5fvaRvX4dd
oHmS2pOFmG2MQhZqTkTjmzXHTj6iuc/Op5ythC8OwyM2vMdpS13cDH2VqXW5u5aKdRLre5lpbDUt
Fh7eErZdV+vugvFJCFKJ7DXo8fFDGtK45EnEzE8hr9oftabaY65ngeuRhCcRoPWvdvkjOcHZdNnU
lz6R8Nwi7xdSY9u5t2tU7sr5SCiFZ3lBXQjp+Nef19EudhONX7LP9GM3vOaVPxN+jN8Pu+bRXv9t
8asTyq+JENCfgsGOs9jNKeqlZmExK6nUiRxH5yjMtkPMee2d8kI4oaqL6JaD08V+tPgoY/2hQO2k
CiBRlue+TDiLPIdn889ck3Lv0530ib8fdYP4pkEWT3JQ0iUCYRP17wIbswxtcM6uk0RI5RrYbQGa
SGjBIWAxthxaBLXpL1z1W+JSkQsYFB2lnrUXF9KJRobXPOBKnFAhjmdF9fu/4K1P17ljfw7FgzwQ
OomRu/hMuLzkwlMNM7iwVS03OE6R39M8uGLMK8dzU3MLKx6ETF7tiZgZlADP7nArfUoN5Mu30BOg
9n4LBI6YvK2ntKA1k6zM/oXQgJph5cTRdhhZeeeL4Ak6k7xwqRh8RZ8bhvcajwH/EmeTOz+kcrQV
45UglOT4mM4gRHufseLpoK3c/lRsMnmqdv9OhhXaMcI7AQzOA2eJGzJAIZYRr3LFNRC2pkxU2A4k
LjeZVuBiGdNOz0drHmaegOtXyAa9oMMevFxs1j5sedd4GFgq0PqOFUCi5Ql8BUFxO8sst2CSVQPT
LqWU9svheoVUBS/64lNOD8zPjaTsVwnPN7Wn52P8rLxo7BXKmqgKvKlCzENt+5s37NVL5REmRrc9
qbJYiY+UpPPDsLNzubooBuCVtgs4PyzlKA9E4DNYonPufbk+OrnK2FYZT64+dDWEqfFBthm8PUxW
mya8/V7SkLuobZy17F6U7lgbbc5KitH72mx3Jwcw8pl+wPQoprSs8vGps875oihjgz/M3jdQY/Pw
QlanGKPcq6syDpEMuyWJhvrQFEWs1N2+Qg3rCxdcExkclT5zf/8jQlx9p8yEar9z5oNlwP/ve7qV
vP0Pf/f0NYX5DfA9RHev7JWqLfuO9uibEv7MXi2CgoSqW2R7xCqgfmxQVjer38Z7ZjIXreTw3MrL
PLb0KRpW9mop330kpUJU4zwuNf5616k6v5uwhUir2pGaeVvcWwnzVAxjSlv2KCzO91XmEf/Z9z1L
Rij+uFDh6lPzM30HwjGa0Z2XogLOfQ16sJtzmZ3Rp/nvL7f5PoOZMk4ZbWjB+Q55Gljk8mBHdvZE
hmu7U1HKc5V5tMo6yEFXAYC5Qcu7kq51QrK6bXJiWRRNqW6FuaDDaLtX0fm8WpWQEXOCei7yeneT
JCNj+eRadD3wdIQaYhES1Tp0+L7hQ9zCNZfwbT5eJdw2RkExJaG2TNEeFF80Cy/DUtnwRHjypU1X
PEY8eQTxC/DR7wGCaoyaQwF0KSdXSql8IJtlFIaYsTvEYtamneV5p8jYa+HVNcawoF4Lhj65eXff
tx/ETBJ9O90HVCbbNgG7C1FmavdSspYFLynyOysH+kksP3Nt0eP6vu2XQyQ90PdToTDsxJ2+HToC
T/Xbc1hx4CUL38lFBHK/UzfMsFaIUeIVzJRIG3nOBe74HmNcogiwrSbQq7rkY2x7IMNG9pCT9xPE
ZeIFr2vhjn8pOc/zc+73o+GemHYw4DLdndnvBsdIP++mIOxFJE3fYVpmDwj5kNoSYoGmnzGdVIlT
nMkCQI3rf0A/qWdaKxVURcn/e+6anyXHXbB41w5e6vsbH/akbyooqU3kno9DaUng0SaV1/YawXPb
UfxOPLggGqq7pwkVmuFcWFI6hTCnrALB8ytZNryhhf7GkKb0S2v9G5o3v+RIeDZ4YoEvCACf/gaN
K2tlX873myadC/hIO5zNk+7e0x5M2NwcGGYV8LSZyAFgsEGXXRlPMUs1mgEgxjmTJOiGSy3XB8g1
+ENDFqQh5RgZOlXlvESP9QRzKgs53wG1QNzIOlf+sr/IyTealMFVPWyz7se1q0bQyK5KdXuIsn6a
hQ/FktQ0l6aVMvpR7yLaDVxh1AQHPiTzci2KGjnEmtE3HBvcnLuWzn01difZTgOb3HrByJr01dV+
gUwMDn4+TGtOcANFtJ440GHdmzA/eCe/QJy18TaiGDjuldRXRdJU8jK58bgajJAAqqlS5D3uyAz2
E5kg7Ds0pAyuqVfBIFVJSd6ymvzQeiJ+xA/DPPTrXoO1+ARU0mDsPmjHGZB+Es4fISTmiXqtIO8g
K4Rp2bUL0fBM8NNInjvmybmviziVFkgcKfRvRPx4y55hqdVKb931AXYb5Lyz1JYboqPpOUbDQf8J
OZ5h4wFbBhagAHIqhw9qeUM5y+WB/AVhJmQUhLoJ4zTswLC1Q1YmWLm7PDZq/0OvunbnY21vD1QR
iF8LmXjHQoeZjZo//jdmEdA4CylZ6CYXDzS2B3ydEW+JA65STSPmrunL/0mqZC0muI7YMyz/qp5j
kL8gVDfIH6H21zpp4xm7aLrFJ+aawbKLdRysFe8QvT3w2fwRgYDvmVWfz8HpYyaBcbVmIOi28KMK
tNk/vzG5qW2y53z0CM+pRxoXWjcPpq6HseRWJGtm8lFepEJ/GgY/mb1Y4MTMphktPe1JpySixV6Y
yoenGkNoJHZWR3mxS869EgjYyAgjPdpu+CUlLZMjixBbPz50jQEetWNP7Ty42Sk299tbVwZNYSvI
Y38xdufdDHkEL15LF2qLRiuOMC70AJ9EVxpGdYuNH3UENMAtPaOSb7Y2NmC9NrYM7rEfQ0DXkm9d
rx8Prhw953KnXX02YFZag+ulIMBJXxTrgMl4K91+LV4IFuiHjFFOytG/vmU7QaKs8V93uiAot+vk
2uYEv8aCfyo5rQK3fZCWETzh41OJG02cW5r44X+nQOpSaWMBTicPzLCPaXuc/ZorzBZLX38qh3tk
oYEUBmUy+Kn6/AY/rDsCf4gkt2WD7kTnBO3/lu1CHq4tMuWpMtIJCbKsitP6u7bcpJ/U76bt2uxF
aX1zW9lCQFWHgZ/8/XpXDQg31Y8/AVc+lq/OOjyecehHK/nyaDTz9QzX50qlJvySQFjmLnvpKajY
xCYNPje9ZfbRQFxfmyoF6jg7OEH1SwpGJ61oyRdzG4pVb0ruswLIfMjQbBI1j5AyIhuGfve3btGK
fexTGgtdBqK14RLDu7AEGzAF0KeEzoE6hqm1+sroFQyPwf+/qY4WfH5hwITUyW9U8k0TYI5LWzwl
t/OticZ6z1BNcdF7VLd4EZfVG96M2R1XNv6jattMnTf44sgndYVUZJI+veemkFFrzVIO58NhKztg
fO180OoT6Frt6XhSkfbahAfbhv40KNWwrDaCVyUWJ1bPUKSLLeUvZhIkLuZ7MVIJy4w3E+5tdkIu
6Y+WH3RvYtfNhIABAsaV3zE+6irVVL/x9yNmzQtz0h2aaPSQAiLwh/UaNM5QATrLeU/lhq/TiSFc
8e+me6C7yueUCZ+CQuNpvRmFlDTAtTBFkBllhJ7qYzmGdBknA8UoD4hZeMmAH3Txm4/1kUXUyQnD
ji7dKOZvU531cQKs/07hX/9wrf5lHXctYfTIFuZK6cl7JhGR4nz5vTYOQEeEDNw9tSLorYNkya2n
fRZw4CjEARobIdaPIO5LE3TvuiVxWTmplH3iFVwEP7JjxqapDjpmIUpR+y0FdGaH79b2d5ZMynJN
5vV5Dxr09AMX2b/OC3G5C3SaCsIXm79VA9iOFUXJ+S3zsEPrZ8pkjOIn6dl+gg2UMXipIQchaySA
Hl0PaIVu69LJqgoLfdBUAWhN3UJkMS5vTp+XgSCwoWjkthiStxT+vFq89ES2Ft/ubDcf9mZg54Ws
KWbRWpW6iFYU6Unl1bUI9DhaInCUMXm12BvBJNG9uo+AL2FNH5lBYYpA+um8p8etyW2KzK1KD58m
NcnE0EFfXHPlDI2CeONVgap7N0SVxgP++NPT0QPx/xLMEj9JuIDE7lyDodH9489ckiAij/xwLSKo
RtfnvXVNoaaRMo0eCiFLLTYfwQ5kKEKqGw2zJhLmyVnGJL4EGZI4dtRC26WblW0xMJ49eLhBojS2
nMMbC/FoC1knDBs/MvZ6/kpC1FukYsCi26EY51gUlQJRhhcehEfA3SG3phHpnP4sOgGA97eXMFgJ
CcvljKrN4W3afXdrcH8X3FUk+M///uRaWwS4bUaZ+Qa4tjzz4sfQC/7pesymApVxl4n6WFLHTC3R
F7L9toXBrTOyaChiea8J4wc1Kn4IYF+zSaIdXWc/lNp/uxlzl67YsaTbI+2TO6Z1Gwt2Cg7EpS1v
S2xQ8CGXiRahBhV04P/Kx1pHni7r5TM8J5Sh81U8Ic+H59FXmmH1gbSqDvb8yAxd7zq9M70STpkN
oPDsTckY4aytNshOsaz4sGVZKgJQy/SjzFj+FtTKFWlIuK+sw0KIKK/kzfiIpmmHfhzfKYewNwxa
w5iaNFvlmO83xHXVSU40F5agX6ICrZEHRm0JKRhHRthZ7J5UWFMwCdO13aEMLbO0aozrYMP3Sysj
9amoC+sFrf8G/DL9g86hEzSnAoZ58bdouTYzSJJMTpV3DmoNCaBX6kmcVxfunUU/4UK03xt/RxTS
BoEct37+gzkmW0v/MGmUHlqxQyJVFGIUNPP6kJR5hNDj8vRfYdGMmwrNmexRxomG+oycdM5bzAkm
u15m3U3NidaXXlUParKAcjTCRe5Wd6dbuf7OoO/ik+BQQKG0mvVUuw8oGoTU4vMGVMG36CC8m9ul
2Ki9hCSdeQRgMUmLgzg2kCGrvhOYx02KCo4Jg3JqjsK9ZXSU8/e5M8DGXhzHIVLZNmyPXa6iiYGa
wTH48SQR9vup1Bgb5iidMt+sUzstmhKM7L4HdK0A40AWmEGowaoMXYYWbayDeFuK9xB+ko1FAOHa
CrRACd3rY4Cc56x0lTto9iIINKNFPYEgj4lkXfxvBGrAqFQnthSn8jwOnQ1ZQZDYcUcuosdE62X6
OJywtZ5SbuIWsBXQjnKUDoA+8yBBa/mqeapkpNvgz6QdGaWh0J8P0Yg2ltNjWKAoVlsDNqBjNotk
QHnSrCoK6BZVxbV5kI4nmW4oTIG4tJRO878+xqWHjaE/nHGO7XGuuEytX0zeL18fEtMl5jBfBFx2
iizbT6Ur0qZK/izIU+HG8ODhIkoN5/rbEjPKAfTS3YLY1MN6RftGBUHf25XE5OoKsf0s/l4n1E6S
OkC5e3ygI117EckBfCEXfdO+Svgs+YpGpiIYajOiZ0ffY0zYKwHohRHH7Dv7mTiblzTQNV3azMdo
rSVr+OYwAwIg6ghUZivZLgwbbP4c38zwUN9aG0WRN4nOa0/fX/nvZRw2qv8KTDZeDO2b9WCGGw3L
cREEfZ3eUk2LmbCoRl7wYjzHy8ZWLwLanaBZNJOHyqhEXoor4XbidraFwCenOelp8LW7YZAmSAaf
9BVgZSrZHUpY8PsoyKpCDYCHnU7jAU2Im4021my9wHREMkURTdw7sBNN6pMs5QsyQW8zJaYRa3Yb
Xf+jkCSRJ+9aCAMvl1v4BP4gWtydyzgJQ24oR6xDPeoqck4MASvFWu5OusgXeOkE0g4BEYDrqegB
fUmjlYhf8EJWU1PmMX6wKpwiM3wmdxqwJ6oZLwX9E9QK5fZHN8hKhk8e2I+Rj+dchTUHX6gx4MAe
wd2SBrBPk1iFOZM1G9uqGxE7ZC/Quewnz8k4Zw6bfIlXR9XhHEHS8UoPHYEm3/xGJ4zx+6FIXlmJ
osAdWilhIRGr6phPa5djFymowvOCIca+umdX0OzKoDjoz7axzYJsHRBw86lTArHQBfHJ2fmxoOW+
DitdHvc6kIgtvJaCob+nNrzbPdgo9/TPY0yGTuIdDUHpsTfHn3jUDvGVH41Nw184+lYn6rSxtP+V
tiVkxk0cZAcTIBt8IDDd5ypTzAmmiHSxy1zZE1NQ58wX1gESKM/W9dlD1HNOHdn/FL8ZrpqYG81d
xihlriKGwVTc+qf/h8+KZWaSJ79O2UYLiHSs1CHu+XQsaHNd5xvfCsYhjFs6tnLMddjuc1KqzkO9
UgWqXNCj1R/lp79aynFiDFpOMT2giUt8BmEdMgrdMRKrsY8GqODCYFJAgS1pJOLm07dM+SMX4xVD
lN6rSQkkeANxZ3mkv5hDkQtRIvbyTvfsRWl+w+vdI/jqohx33G1zqGN5gRxOwZ4LjgW0KYzeDpww
C4hwD8zCEIsY2NQETza2oPnAhTKAm3EVuEgycB8fbeYn2x2fn0JYSsRqz9I0Y2sT/wWI4PBKv/I3
QcJ0k6ULxAgXntTZSAE9gL5x1mTL6sxO7bCtPHXIRow9ziyld8nj/IBrW4o5jzxwZX4v6+LY5gcf
ozhR8xsynXldLzLCrys3fH74m66UATUq8TA+K+hYcgzFL6oBQ4d7ZH3QkXdi4rs0+F2aT3iJf/Xj
BnzkPxEZssHrBY2DbMdzOJ4i1QLaDE/xDuhsTwWH88pKc933rmSkgWAMXhuMAXb6pFi2xiThLJsV
/IjM/8jv7I8ZhZOuQINkxqzRub/SJvqoj/wESfF+dpy9atsZ1MC5n50WpI3I3p/IUOOJjUALhzSS
u3ZD9a+ocxEo4dYVkjPv3aJWFt7NY9goiFxVNepPOAUazZBDrxja1YVg7hJpzyouQerOJBrDP5BS
rjHhcXBk+uhAF1bTTb72JeoYb4f708PFw6vk+lfofLFSo1eiwEHL1uXyHLN6+bWr/MLuxEugJ+dq
VxjqZ7wWbtx6Z4EDyFjWOHqy0jU1kSyVW8b4eYgtKdEOxEsMR3r+WdImF0+xLsaFrKovOfLvcGEv
TUOh273P/R9IQbGaIb+SpW4/w1wCWn42uZ5ZT7KpdMmszkXP2ws7HLF3N2ekNBzVbcU/na5UuE2a
pyzolsRmAdGLqA7Y8n2zP29YHidDJzgb92Q9u0WhnwGE8k+hTL57CEbCTckltfC6qNAHM2cZt54M
mbxINXn/HiorLlZypDZAGDxK+gNLC7em29K8rXamnvlQMOERUBPzgDafi2mzFKzrOAZSJxmZ5SbP
E/P1T0FKGIltbtn+Ti/HphnwwdUHXwDajh4M9c20GkLevJlLK20OiMVv1PWwxa3HybHAzWwHajsy
RfBWy3YSkgz/SyXmVHgRe0pCK1bHMSI/TYu6sjpYVQjo6RkwtVXVP4sYSoAopn7mNwkIGr8rcXo0
gSijcrCCIz7Q3e480vGhrF7zWyug+VSRUQ0M4gXp1d9RPU6XpJyVLCS+oZN0h+2GvDdqTAJYnY4A
N+kpq9qC72nm0sB2bGnwj7ZGvp8u8W7I7mg8VqHbt2iUoUcNsHux7kC4P0FUn1PzEZW7cyV8D0Uc
rkbf9nHWerOqhgHdqor+kxdDtpbYdRA0UaXZXz2YhH6MiN/Y2pyM8LN1XrEI8KGp7qy6LtbHE8K5
4Tazeg/883jg1w1TF9ztJUoaFGLWo24XaBxHfSVE0NzLwuhjyVZJggP4x5SEhoNUL2VU0Z3Ch3/m
crM8UzYpd8zg5l1tWdQPdEylnD0j0s2kMNRsu43T/p429jINnXAxo40W2XzRx4BZ+v23m/AikUw+
bYYrJcEULYYd/51V22KfdvgFcqmeNRNyHwhveqm7K991DnlN5KGRYy7IqjN7pw8Ab4yVGDz7rVxq
8/sO6PQrM00Tv/ARfEXS7TB+0Aiy0lh84j2paBpkXY9p+ThXpST2ywdVU5+1VQaLwo4V1Zx1JwLL
hw7v4FbYLOFAtPNfKTnp77qAqR6K2aKXrVOGzkUiwFQAEEDR07fFgKCarNh33kJO+9hcwtjB6QIP
7MWp7OA+MAygRxL9ruZhH2fQDAqE4nrc6fToPBr5tManeYJl/zJDO6PabTgKVDyECSot8XO08FuI
+X35TliAIX1/rQZ0vM76+dk4bgfpdAEXT/CmA+QFwS4ORUW+fy8KgKDMIiARPV17se5O/V8VgLKl
D1MwvA1OcqdpBGSxaF4aMKDF/SLGlFNrIlspXE9E8BzbB69xd8jSKm+d0Qvu88O3G8xiepETWS9S
qY3nlcIY7XsScZHQes2vSz/5jyT6zWnaNVoYs4Pr2gAt1bn6nSfOHmI1jRi+7hmJb5lY8ZGLhRno
XLoHl+iAKyP1AeCPjiC1TcBz+BGRXaOvS9ZzO0iDGTfORBQZ+ZpMlUrKHaDROjaft2ewqydJZdDB
2q7cLA17AId6zvs0t6OCeERG8jVMiw7XpFaw0SsCbeZSKayk2EGNqwKX5fcThyUHvmk11a9GX5/C
GgXrM0GhWOXx4snhk7nzMki9rzlYNWmYOhRRxJ3/wXe3c43wW8dXOuh1rqsjnvkW3sTl0ylY6RQs
uIg8IWCjm09lKPY5Yko/gA8+RUrYxjIYXb/NNrlL9jbYZIrI+1Qog1m34DOEoQQt7Dnj6IHm8ZGi
gLVxDIxO279O3M/ffzDrfrTYXeJLAD2LdxTjpngZBdvrLsRvDcddxlHUxj+FNIbbsrlUHOP5s0W7
Yxzgr9Sp58cVXiBIaEjKrCLLg/dxAk58+L7WPQSOb6RdE/ohXd6upG2yCv6elrpX0eIU4z8Xk/Xy
QTyb2L6Lx9TwD91+xu9VZt6tc99aDaFe0uF/llcdy1qafCpwcnjju3TVlKbM1Vm7mdT59AdyfN6Q
4J86o0kAM5tAITyezPNgUOIf/OBOLLsq6Hrc70z8u4FTkCyngPDKOY1p+InZNREJ8jC586M72lGJ
X8dOXtKfx3zgy7GdSwXaVS3vbHY1mh4Kz+kJUxQ57hfqKqss//SrwyHzYMujCg5jTYPwWHbeox9B
uyMlxjVmT08rMVqQCVaJNKMuXxnZywY1Jsc2uIBJ7xrLwKBWaYwbgIrUF35JIx/xNkgKWTNNyq6j
uAAeUd0YQLAiFH58ceRHn9LEywEpCYdleUIO/Fi2yrzWvzhjz8dl2xssSiNtdjFZon34FaCF7t75
ALVowKxNXBLqHNrGUi67j54kZCiTX6y1lb188/TgccoQ9NzHMhVH4rw0F7+Qa8gmQokxXZ4v76iD
IpWvCKi+osmDIo/8bw5uMd9uuiVSzyC0l/C/N++xf1mO9Z6IP2hFJ1b8rqD/n0zMR65SlTDarYFd
4B32leX1M0mg8VifdEpEsF4AeUoncuYXRtswqWN7VhSUVMAVY7eE0EJKqJ/pv4kXJu6lvQCJu1RK
duk0fmmX4LN6KEEgIgOvEEeC/V/J/MH391O11a5kIWZxZbR5mVqDvXo0XywdPb8NSSvK4UYBbISx
VKstS+DenWV52+7bRVVXz6Oyhyz7u/5vjRLvljg54aj06j4QwkGnF6tb6/WWFaDIYvQ3OEH+qcrK
93jnKhjksdQtBOTgrf258DrGTWnQWSZ1MH1jX2ad06XronJt0pO3TYhoxevNYF8K/fFsNu3ToERC
lqRSpF+wwKu2n3UZ6/67TpgkqDMLMNExxSQD6VB0Q7Rp9AXds5RHBITXXR3XsljvQT1IhWx/cM34
gmP6Do/tBu4stn3aIjSctlKLHbAEqwTR8SIMmZ5wvnWSTJPWxjPTCoTbmH6oNRX2mY0cbY8N3XYG
83KfTt+gaPnkFc71V7CYuW4rxrKzFLnR/e9DteID7HxtMce24f7E82Wy5zQ20FNAxPuopD0CmNZk
GsVWFyZufRegy1BwKgx+ePevNvvVchQcWt6E9b+vO7WBBw0yb87HdpRCOYFKTWSC5NF/GEZgdx0g
ajCxzVKgWgoPpdiwtdC9N1+S2E+eDyVlB8eU9eAvgtCSN3PKOgCETy8k76nOeUbYSPzyJMiTTHFF
cFDMUc68347h6oRhexrO5evJS6Y/rs0kndpD1J3/EYcKMikn2mVISKAYd0uym4r1nfQ20zlIefX6
hTh25EaJOCjMMAeg8NZiKoIB01SOhbsJZ313QObHRcGunGBkKO87kPgIDJHjAgm83+sJukrGmvyt
8CK0PDnkr7iK8cHB8WHIdFTC6paqoKxEyvAd6zlWpUiwdlZjKg8wgpTZB9LR1VRfZZc+KK6QcjnS
zKLpPP4BrsctOa14eCJ3WRLcKDNHdYAD6arf1H57gtwYyOjB3pl2jFIzADBhiw7B18eycW45ZZv6
jztG1wGtuZXcKAmqIKFesbQEG31AUP8xuw93tNR0Niq3K+qACrCfnJeFAJjsICFgPjRjuZOkzaeX
idKNiiQ5uLJVKZt5ghF+lBfp3Q0mj9xqoRo2ekVvaLD4i9dUeYDv47ajdSktriRqApXEb5SaMug4
X+fGfUInCp+MX4YD06byoqGqb2B28SsoMC11PzhWRLCcOoJR3yoK1X99aZJvAtOQCKGZeFGMFjku
34cvITiOn3Sa2Zdugzys0PQSy4LV883fvdWFzTjJIVzC9LHFvPOsGfOW9Ry7frg1TWZlvOgse+q3
+t8lFg1iJzsRd3taqnOI4aA7bw5j82fmiA12KHroWmQ1oMEHEPZ2lrGVW2kcUg1EwLhQCIrZ7gDZ
leDQpr/2WSLpBKZjK18qsTTgLGnwfW4MKBqKxc8cYnXkPZckWQTku8LEul0hPR7vBnJCJFxkA438
guAOUrcLcAmjwB45I+aHaGKqOWKTkJPaI1XjRevvcuXDMKDuF+BPlHyYewQLtUS/4oKSWIHjexfm
7cTGNkh1U/syvd1tpwgSrs6rIJgbUabCj/FqQRXgBPNwLg4UP/SDunDDi4OTu/RVx/3N/jFw5Xoi
049aXrTaVvvaNNBQs/NX9qsw40HnJPB/Mrc4+/hsFalRMUc7yilmii+i7ldveuwiYvlrtzCdVmJZ
Bkc/YYSiNOLF25PU3iWW5l+6f3sq0tCFU0ysIXFtalkGbhw7LWAT38DoQ+GuK3mR4ncN4UDXCO90
YSnkZIFmVMt8zNGOZd6S6U1+592h+y/Tm/hahh0UFpGgmD26jYFnt7X1dqi3cj4JktYh1nkDf/vL
ATFvxl43rfxcmXaDXiQjhgMNaxhFLVmza33KlwcXUhxQ6/pqEKiDQiAieQLVQqFWiEl1iItkttxn
5Q/LJTbmUQW2WPVO6FB0ULj7hriWM2QGViM6AYvvGapHG5KBqCyIOT5uwBgr6RiCrCjV14shZnyS
vJT2/FW/5GM2Iampr46uHXG+q1k7yCk0ZhT89HNSrWJzzLhh/fQTn4YwPEC8mAWh6REINlyDiIYZ
uNHo81PR1Dp558Dg1kSQJmeCZarul6NtYlu/Kvx9NukkHxjhfzp+ekEwz21dASJP8tOXL6hgPi9i
2SLtDm7UtAciP5GURvV4iiQ6aXWWkPQMEsAWbaa256y0mbYvqF3YP4klVo8pHzAu/GMQrtdaYvV5
MHEGaWYoCoaXOO489+p6RScp1Ykq+O/XLILDe2Pd/HLb4cKgg3Ui0tunQAKnTY74/Rp3RDfivPHV
DFA8AKAMufFIQlJu2IRCMM36PjqL/LiMXBeFaz2i2OnmKTKdD1T3HJfQeubRUOdQ+cyJcEdjJzkw
ITwxf03MEZi95R7jx/iTY/v4atfw98rR1aoT1jxMIVNsach16BpOvgAL7+HOjvQFz7KvfVYmr55n
I8Ysr5sevsO75CZafGye5c2n4YuF+Kpb2mT6QoBQP0oMPDeDPojbuKUaeujdqDlHOOzwXcjjh4Vg
EqI6hTWWsus1lyS431Y5Q9MrHus1i8E6ivO7u/yhwzVRZJc5MlcbTnTp2nyE5Ej0tZ9j1p7hEjer
txHVLrxYfe1fwi5PkwlHXv2qbiyCpuqrB+4SyQ3xAI84Fqv90gh3J8gaXJ726/RJwb9WZCGxGT2x
VIgBxYpFf/m2lPfTKff6CcEz7vIJJkTMmhXGeVlICZapwdTrObXC1yXdjaIUliq/ZpAfNjOgNW4v
hF330ZeKK6YMDmdnMNXT1MC1Qi8hds1bOD2JEYylqklDWGDFAygaB7VBqT/bIIHvx0Q4LRr1sHkt
XjghWOapGuxDiwEygsHcjEtuFAJcG4mQeBxzU0moZth1YmcapDlqmfCsl8l6jE8LYeVBwuQLAZFN
Z66L8RXF5DwM7WiaSfS2ip8xA0Smstg/v1eMub99FhyrTvEZNqP/ueuj/JlrKCT+DVRJ+mp6272I
Lw8DcNqDEmkNpBpd2gf1p6ooQE+uvP8KyMhj/jhaMiPkAoTqWzQOuXCSgqYjzc234EGBkV6GXT3w
qomgpWVknxaS//OiBTV6IClnFiMo2mXGWNUYsBPerRNY+VYLaCbXONoLRqbTLXjr+4vFdVHADafj
0Jmrfohs6JVELwA7/H15LyO/V6B8sAYKuSCKNhI7BxLSaGu5qJOVcb2u8AsXhC8CSArhQAYicqTg
v3VJgBMXv/zbUaDsvdyT63LpESp2yMzkb27aBxa6i4wWqnARuHbL5xwhC8IlU9BaTqpAqkjJIAge
6u7Hx0bdsFIZm9LBBJPqUhrVDowSJoLatf0/gvGzu41cSuEHAoFO2MWBCEsvwOUkok3sbBARWpyO
IQrBVglXrzd0raQoOBUzoo/Q5JCbzEwV4nxBwy5i7JR6tmRbHfs5MtMJN6wlAu60L+87m+vq27Gp
rVgJzx/sba0hBwWw5cqZnhMy0pG6X3QsmZ39yidgabtOxajGbs44x/XxhLSufB4RmT02ve8kOlN9
dNifWVe1rs46j1G/sQNNL2cf+tP0I0BSsMufEzKc79rm/dXguxN9E4QDyeJbbn3Vl1d/4gs43vFB
nt0FlHz1yG8uo/Yk90KU9LYmgAUpzizLQnK19E5yqBuYGAu8FXLjpaMHeUTOGXhEkDDGQKv/6jot
wCENI9pQLjAOPLIr9EPzhWCXwBD0YkUf1EAyBJKVg5auHGGJQV/xGNpW2jS36gX1klUNaI5yrN0s
FJifGjeO5J2uBGSqlX+/dF4Zl0PQws51OTsKdRta4TpwS1xmSWqy22wjdPEYo5yn42XngXwbYKHw
HRb0+uvEJts+qJSb3+rqf6Ka5CR7wM8wk2nKoyV24IiBB1Oe59vTxMoPCSG1Oo9gd1yKLJQAdAtT
fm+XDHk2JvLIcV6XtA77SqyY0ivV4aTnD5FgZIn5voUGz2a/lhEbQEerhUCah9Skf4+g2XmCaNYB
DBv3anRlvH/RJeaHXkGpXwQajw34YjTzIdGsy1B6ZzjfvHYiwKqfbY9QAcZ4cq23K3P8DTAO5HMM
ddRuFeHC5sECijl+gSm1A3ogvQkHL3Jeo7MgrCs8wBmxR0uQUDHMbVjTGx+x/+IUSGkewcJDG+P5
iqI/5KWa18LxSaqBw30X+4Ygv9AYYxT2nJkDFiEHR13FgBfeA54Laluvx2aO+2vQAVFrg81s8Wp1
EHIUAqu3CyDSPFF0a7tE/CIrGO0KOsz1Tt6iKLgzc9mDMkI5UwDlp33Pc1NSROfDAT87OX3u7GwQ
8tpEUzicfM8Jih32ImJlHr4cdxKmV6W0gc5CN42SmSwKDazrZVnSPK8l0z8FOr7Nt9zZ4tZoGm9i
77B0pa7yEqHysGA4BfR0lIVTAe7NSkyndh0ojH0luN9r9rg0xDcIONCshAUFrbRk6Bua6lDlJ3hY
xdOPZkTsDOoYSfMHCtWh62vCJdD+sbwbP9ugNBfiQbECpuzqP3Tf5Bdbd1RSTclWpYdyzv3+/srP
XJfJqLscYbXDHXv80MT0D4a9/OIBE6AcHI6tToKLRN4MVg3o/YtHJsBESprix2xhRDapMM9RqSps
uy7/0oTpyam0KHqMqmV9qND9B76FapIZw51d/9Dj+bdAuhQY4CiYCxfarWukXuTK7h8iNJ2k99TV
tp/BpjI3DBcgAAzYO7BQQX5CdLkDPr5yWpHyIz3V436oOu/asNip9tW3UIM0sRNlvMzm7+lSn3eE
4ysx+rOZqmwgLwFsVUHPTONTzX5McnNw91J0Sz9xvzZlTEg6yOjTlEKGqh9iXR83a0/Ld/8S3Gg/
OIIeRKr1dg0k8/xYh2TVLqsOqZ7r0yRCKjmFeDWoUu18y5g2lwI/Qrb4HJlBqCqUUmFiTCOwu2HL
wuOFFLVgqw5vylvv89g6a7vblUS3w+tlV7kGfLBYkJwCxGfEp1V6ZQMt8QMD7Y9rzhLRZk+1N0FC
F9Dr/j1E9Zs8c+qCj3FWfcjWJWm8xlygz8Mm+Q4AhnTaBy78p4mocWyqe3HEVY/jHHR+f54gxPNs
CixjCPsFz+yeyfok0SX6DezLoaqPf72snRdqo3lcmNHudrxGBfM0/vKJwXAsch2mkk6iZRMXrCz8
X+WXqUH2x0VrCp7qtJYAnmSCVyaY23A1oqn1rDrDuXD/Tm50zJbPw8X+wksDKTgH9wSxYiKjoqDk
xJtSWGqMsvkxqyCJ34tom1VoziPWRS5V3I55BUfA8dP2wSkK0q5KVWI8aXH0Ov7ucpJR6+yZqbQR
n0ffCXHVPN+GVbj7wIeAscgAOB07b71XT3bV34R4e+PoTZPz6rT6hivaAJzpwqu9EHP1rOJ16k0h
jA2b+BCy/4uIE2RdT4dBymVRavjzY1g2h22g4RtLdoKsxDrcYGmaCcR03/lMwh5PzaYW/HTdzDF8
//d/xDxVxACjaPiEVaf6d63GHhHpHTHckqxPNnpINHt7DW0vP65v3bOOYMHyoV8uAkqKXoue/mhQ
h9eZaoc0ndb4xnWaFwaOw1XqNKth9RyxouR+3H8npfgvArQRC+7AF/oKjPZg9bcetzqYtOi31ZQv
s+Q4hFS7llr2RgJLWtsNjZKAB9WvbqUclUPH6fM8iJU6kxMTBKEbAWOzgTey4vO9C4pLQCSzcLso
d8NgmLBgzHPSGTOD89Bunww2KI7Ib1Q3dJjyBvu8fnY6P3Mvl6P0Q5cb4a5r9c6/WMxBC48udRcB
+bAR4B6iIkFYesT4O6V2S5NAy4EGXgBkJuoYxyxkiRA4GUTHfogZFGHqgP5+t2rmTMfsBbQn6u3Z
ZxGsvRoDUOcXase0TIDvNUb+7UMS/eqJuASp+V3Ht5ZL7e3O24kWldPm5MparU8HSUYnHZf3isyN
bri6P/sqANHiGRd3x9p6XXTdoJcKxkXHgrIvacs27Yie5EYH9hijxrogVywt+d02K/rGeS6GLZjK
QT/NyyN6XBM2Llf+BDMoe5YOuaGLxGZYU4+JWQWe666mTAoQR21Lakn09DRfKrTnJzSxbKAaJ19v
v+hG2a/ct9tOds2P0JFhiV6gE8atam6W9sDPz99x6cWliMJ+UUEHPQKlHfUI0kCPEX7f2u8eh4z1
VNMgU1bwWsos2b3vY/cLUVncLOnsPFwuAhbbgIZunqtbXnz3WPGrXrpXVKAKq11fLdHf9JR4uPUt
czUjKBCw96Lo4u46PxtdeGt+kF0DU7kfE5bEvLTo3a3WD00h6eY+uyO4Is+HjGo31CRbuNYqIBsT
sftQmFqpFkVdwf6doV0dDzvFpyBVIAj3PVpbXUFCOm6k7LsBLxgdi07IUNQQIcQk0MdM8pyQr/yY
1VuZET4286ic1qdIErhr5fBaOyZvgFpGvhRhoWUV46WH0YPYIY5VNIV/6k36qoquOOsTHJvGEOmv
ba0rQYDy9euuNek/2LQJV/Dk/a6W1f/oq/Nf5CIT7soLd3qcLHJbET/w+5cF18+mOyVP8WtkR8UI
/ZFHYUgauCbYjWv6OZmSVo9yaklu9fTDR90chjBI2Hub3V6MNST+bVvvSgV9d2Z3XRiPbh+Fra0V
/tSpT7H+MT1XVG7NI5dbavnc7fIPEfxSCj0lRlhh7Y9OQn5Q/+wOSZszJb0EobD1nH5AoBxijMou
A7UuWmMlC1m9ZlA/Lf6oXUBOLxjrEJEakNqMS0ZOvYeBenEcOdy+Wo9i2cGN3qwpx+8q0MAHddu6
2iRqw4aXMkaSXKc/hMfD01+eSyk+QMMSBT3pUYFa5B8JgVWfKKIqILaL4Ia4AywL54p55oxhGRG8
Rb4LtbvwQdb7pV4zA3ONSaYH2QZMUe+tkt0JqwnDBG4P6TwcgCWiPxLC3faQNqxV6gOanFTnzy9M
VuUdNTPGgn+AYRJyfhBeI4kS+pAgAy8WdmDhi7PMpmtxK+TFh8XesyOUbFf+5/vwYdKlh1JEgCEo
+ti5NjtN1AKnhNnkxEPPPl5Hj8ueYBH83ydmT9QZ9NU1HPMcBiDLbUmiJFpeVyjkPfhAyQhFFfLT
WLqgflgeiXEGZcPGu7AnjUFmN2ZmIdIcRbig/zBLL+Yhro+Nyf9YjO2F5cJFFU+iLha8lgD1vDui
JcG35bjl3uAlZhU/PHrV2VHpQYPARyddXx3RSBmQ1Xg8UVaygjgmHYQGe4eKgV2sM9xB5PGF9tPf
W2ipTEzJ/5/pnKZy1pWkG4p+hWuqdDzYm74N2U01quyvbbq9LcY0e4YGdBwiSHsVIE4VJ5WI6wXs
5so84MNt/8LGLjljlxMM/GH4uJtVMBZMqrjiuiRe4dlB0knThXWzvO+mahtFPlh0heq1Fh5/3s/X
SomUL2IVu66V7lp5qcwVbl67fhjUiKeQ4c4TX1G6tbOr++KmbHD0d55G+7ossKUAUyXF1Yf+0ZX6
gMIsD+c5bFqOiXq9L3RfdL01ZLxLOPvxPto39lGFWLGhVw1ONi41gQj+S6TQFEpB87wDgV77bcGX
qFryF8G436swhDr0PL06ZXLDU1MrQdsGjxzTdr1BEi8tko/oYHNAIDxnUezkVO1B+xW9FvA7R21S
avRH0RaXrZbMYF8YtpFPGT+RdYFxRnpFh1nOMBgDpOKmqSUhD/vQ8SOvjealBMoDVTP1Mxixiew1
3eAg5OHiD0XrEVVgXooz7aoD457TLXD6msROiI/v0qYnm/lT9AfEV756a/Qlk5kAqB/f4YhFsY1V
/ax2CZaup4TaNZsUaNuXf3C1+w7euVhDlGcB+6m9ydC1Xe6bv3pUbijLXyZPwvogXhMfFubUlL+J
1X0lV4+4RKiSxQ8Matyra6wv1pFTYd2UQzv/iOAFaoOQvHSuwJc3KgVDmL+RbYRC+CyOd8YvOqGe
PvuP9MrcwbmVq9qbBpLEZpUdtKnQgyPzX4YpuPaCzPVPTM5ppLZj9z+VZb9EWRBgCcr5mt+zb20T
8Ixdz+Oqu/sI25LZt9b6gGeTJxlCfcn/8dMQCfXzwca3P/fjGaEQMhkvdpVibSTisbngMe464O7g
Ln//6NilkdofakRz9etZ4nI5Oj2PJXEVEaAZ0aC2yhGw1PCFA9jEaQip7AB/St4VrhjzHeh1Dixi
FQB3JbDCI8daxifg+S99yML0WLWNZ+yuCSPhlAq7Ckopz6qC1BXnCI95L0Hsb8OU9/sxAhlzuy9c
V98DE36PbYKe7uf3LIFacx3fAanb60NVynKXSDJqeV+JEMXL1BXJpmqrSlqrp4P6DVmfTgE40dUq
02IFINYu1DPpq8CKqWbGAnr3a3iMfDEthzEMnZc8KstrbCo3s2fYDxXLs3eUgy4b6TFd/jl2pU9x
uPkpLktT76d6YwkU9Z6QL2vWUc974WSZ1jgHv0C+yAYwuB6p1iGKWJ6FGYpuislsc1LF39imgjM4
CnnoRNMg+d8jqNs74wPhi5w/Opg7bEJbnoVIf0xalfgqksR2NMP4MOcpJMrPZl6DsGPTg1XXbt0R
UXQYe0Sq1SUPWE0dp7deBxgZ/1ecwKMrdKadIQf+bhJsUHehPxFF2vUu+hx3YWk/XEftbW1YSGWp
M26f+Am0rvqpamzet7XYMuaGyopNKvtncy04OtNW5HAKt+Xmnix3tnCzx7MPON/Dqd8H+tAizyEs
dgT1K//nuAsPvaPe3BhMqSjSDQoBDTwuv0/PcHRgKuerw2kEwLJTwyNXdRijDGMR7hDbyoeHvJWP
j5+LUo92Q5g7he+MmGSDXPsWmSuq685Ulm20ezJVHR7y3BXuXLj4anKWArS3kGMN5i/5X46tUf2h
/OpNl4kr9v5nRDR7HeRLOX9oz4HLo2WhAsFF6e9Vdg3HvJ4Mma1WQVJG5m2dSIrTUxXEP5xdTW5q
sWQmP9SRkQJnmiUgJt6rxiCe99uuWOd/aGx7jLXflDnPJHQhNMnEuGJQGKpR9zdS1suv+ap8Z3di
Fb1rZ0YpH4f5njbybA/MDJzr7xya/hD6NZRPhGB+i4/6c+ZP3xCEC7qCQiSphHEhqmueUEQs3Pn3
pDaxRX+nm8fpYnX0POmPWZZkgnupMx8ttjkdvKCo6Xgvb/j0XiDnmc6KTlZ3dKhnp68ZFVjJ+Qlo
k/d5mFv/J5QUjU2a5bFyKpEASSWxOAK+1mMjywj2gA2XZMAOCsKvtaVu6426dGulwjuS3Q2VUZaw
6ADmBpdvfpqgY/pEVizFfyLRZ2MtlLJOLqeZUY+z73SHL1YDrBU0COABR34HT9llUcKSntTNzwVM
UhP5dDegbdcFdYJh8F87ZPpxpjMq/FFXxKvlvVhrpaARK8EMFYoHIwtstbN/dNVj5iAF+d2d2YXj
HEvW8cgzx4COmW9iOjZKeDmAsVtN3+tafuvjo3HoEk4HaPBGjOgq4V73otnEGC7iuuh9x2XaVG83
3eauhGe87BOFTCjK2iNlPl9AjB+C8m2Z8/7JxxW9wdS34/HKrIQ3v4b4DDZuDPL4LxaVI845ah1A
rLKzQA2VjBLLsmHFhHhufGIxDQ/3hFgj0s5B9tKuZmCJGVYtuLtkYNVqyjuvEFksfKTtKheC93BR
z04/HsQigh2ccLX86M5NIOjV4+sX5Hdv3q5Cbz+nr+5lBByWSU+J89KijHGa3MjYb8c+A76Qd3R2
UD1xwFnZhWfpB8u4p39soD8tf1iGjeXiq+BsOPBpjj6D42lqjLPiwUftgs1hUAblTOnAStU3bOuj
dBepXRTIj5kC4s8I++JoZXrNxwgWUnC1f2p1ZuqcOyJeBR4HnMjbRj0kEs0e5KdYIY8+Cjdx+S+e
/s7XbYuda45PQFdDWsy68nEKqD/s3I4PRtaN0FBuOSlgSt188TgYF3Ox08yL7xqlyBKAGkltUpMH
1BCRTnXRonaI7ngzPyyNiG7itBNu6gGOK9cLxJKVA65Kb3WZCVFV1WIW24EFBEVKRG9PLfA/1kjk
sLJCzKnv1kPgs77IXxAxzAh33pFT07lTlR0pjMACZ0JsCo3UMPcjKkSv+2TGDQGiU77NUAV01/iz
ywxIiZph245SvnToiSn2TgfFa/a0dzt8Rj3ALbVoRM/Twg51I/fzumMmeCcujsFon5fPd0cLMdVU
70+kvzPydiQ689NfzadTOOU7f+SzJmhQc9l7iFRQGMO57c8YGFRIhWYsmwIe7seMJlJHshazNqk3
ozIMgRJVW4/YY4nByN8UG4uvYTF+ik4u3Ts5prNzIoc7+0kbLwfLDHyoGn9/PiIA0TShEadN643T
nI/7b13cN2+Pe8Znk118Oeo8G7EpwasQMieSrehbOWkK0SoaaIqryxjza2m9sYDDGl6ZGYXiFq3O
/UapaugvbS8PnNueZlALqM9uUawLLEzSm41KTCnGycjVzRdCEmHsyjW5T4zzKPcNTuzYHR/k8k5N
myNiZPR3px9BDORz+pZ2OwoXdBkfrZPs693O3tJAjOQ77xGiB12Py/J+jLMKwoFFHx5N3v8gUBSO
K3/EXQb3w9RWMdzQ3xcc7AUI6hVzyEY8lrN8bs9OrjfHCSP30P/742VAsSJwQ8LbC/tVt5DMhyrc
JJTU/vevvOCurNCIsAwqQCoi6qu8ROX3pOcreGB3xPfuwWZ89nN4wOUJNzcXaLJdaFxlPxK4nFTY
9gLsgdIWOGjoJu4QITxaEmNVhfEFdseliL5Toktgp59AXQLgp7V3sVkIJ2olWhbnTVXpUDq4ldl2
UciMYy0LHdiBLN8+PE6bPHiEiG8wM9oQPIUYuMpWALcskdd2rl/TkIygWqr7Kjmv45DrYf+FMkcQ
b7IglGhl4wLx1gVrWj1aLv+cylOLu2VddV9F6/aDlDDE3v8V3g9kj1A/1xukA9NUdUOd3zLn9LC7
qC4J/Qibjdltt774VxJS1SLyctvE2e2ugkfnkcx+caKvqRlHxsFAafokM5T5OdnR12qw6U1dd5n/
x3D0RdKdE07bi0HbNRapZuBFoc5gvJfOXwsYwFhsOLfxPogSPndY967/FXPYl1uNuPLIzgjVePWz
l1QLiiBR+XJwQ/UuGPu3Qjn8+LfECtIqLldxBL2dMsB4BqQ/UyH+3ljZSNfB4zzS+n5I3SVBCWI+
ZjhHTZIr4ckFBrsQwueGjfqgzIr3vABmm6zIfbOklliePoGDstRBsWJS6VkJhdVb1pjl8qkTuE3m
ctsTTsPCZqRqp2923jl4G4gKYVZs+E0qgAJKLm2EXRETwJHt7NPtZMhH9TstjDEA79Iolt3X4t+2
twArzMiePzz1U4qYazeuKWLP/XItNbOcWrfj8Yazv1w4FYouSLdKvapDtvwXxXnSuCspU14OcJB3
/r1Ps4CopsS/0a9X4nM2zhDYuhrmKsnMts8RuEP3W2oTPyIA7/fxs7F+orTgnPa5mIU7XdfkroiM
myNLZqPJAbeGdsTc0zZIS4+OmhTfjVU02QBrgPYdTdq2RYMmmiivwkWccBfTo30oFGDeRl33d8RT
SBLV0IVEsOVPBCcXFSwYy4+CG2038tRjSREjkwFnPf5et7bjgeznCH4ndlWNijez63dfh8Cllkra
ThzKQR4j/ImTEx+9i8vuFiOR9fI6FmTijVqIBGXPxQb3+4R/vq8d3nT7LJq6hQSnH1TbF/Gb532y
TbjYKJPKSp45SPIz6j5j6ukSF/9Dgw2f9hxKJ4Sr++HZ0ojK9NTpQTamYaEcqFnl8GMJt+JT633J
Y69viUHZ+zdtk9kSNwZpsK413zZK9SgZVZC07csjJXpxlagYLVJf8Z9UiKCJZ6yEb0sU4KaZZsBz
wel5gYT+5ArKaSvt6LcY7lIppPPcO4HlaU6lFBsfmCl6gomMxRXeOfckaMSkYC1fniGS0BhY3Plt
wzYjYSTeSzMxWiG74vHjMCOj1IRLlFSFFSfHfre1nrCZADVuCVqHMyJLANbbMaYEM6XEnW1iyvNd
zaw+Te30MabUsQbfJ83nwnqiFIA2iyHpjiqNEiR7ofU4672kO8qgKYCc2Y1qgu15n85JTIHmug5o
QIeG66M7mYzsVqZMbzAxZIeUPFtKuljRVFAHiz038J5CgAJ9tLOXZ8Dr4ahPa0CTHHWaXk2psgIT
FDnjOxrvCu4rjlnp8gjpnuNh/DJMEFSH6AuahsRla+KYHOuzIqPeqLdEx0Uz2S0DCgvP3qU0PoZQ
j/hMxOfbAY65njUeaiPdTMnv85bBimjN1mEHzJ0AfMjEZrXlGt7roNEt132nIyqTs2jLyEOd8qRq
Up6RYtKe++ess/T7KhiH8WvQ+UyeLaprJrAkJZXP7y+e6BLGngHHIEBE6GMACA5XD7OZl/17rl1O
fkhDGYQv8H1kReBDzAnKqnCnfzLN3xVS7f0pMWIdRtMz9FsACFvgdoiDda70S490WBOTOcnHl9k8
KRuBc2tFKsd19RLofLhKOfsaRoptTxfct9ysfxBUDPWJasCq3fCY/ApjVOXXV4570AP2HHc1FeRZ
WcQlJQavY+zkFeXoDwV+RePiUT8iQyIa5qXsVcAUH/i/jEmgJuGbC1EVpOmZFKSrCic11+nETKBm
k5GBkzuTLnFfodryFiFfaRIzDkjruQI=
`protect end_protected
