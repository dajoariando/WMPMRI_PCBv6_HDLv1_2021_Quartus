-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
S0sjO8X/Tz94ORUIlZAMyUMlcSOM0KsoHiUyxHkm2T5CmoLZqfmRaTZocUglPDI9Z/6r6TJ90N8W
SjXwLCySmc7wUHUSA29CRfgLNkRN/qLA+4YlBj9QtU66JiX+Tc7K7u3BGLWr/1sosVHuBrLq/s8+
3SyelzDgl2iIEwSxLpNa6Dbkx3caODJnTHOikalCF9IKu4KzmzvC4/1NGHr2IUrujtYU33+i0Hdr
WbdmDhUTZoZ9neDGvQVWWeiiwuSAL4DNJO449+mAsD6GV8+aQAU+f5jZKdH673LtmlNVjCoN6P7E
kKhpbsgL+sR8r72DThE9/e6LqJFa0wlrs2i9bA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4816)
`protect data_block
pSPOi0zFQe617NQZCGKX4NPtrY6h6hZCYqyvSfeEofeyejOBnLrWw5AtRGySA7+/PEgR2Kkttml2
7jMZMZvGpur9w8mRdFuJ1pdWZqrSaUWsv/Brw8FAvJwtyvR1mNuBDGBtPucftBK+CDVbmxFnclSU
IDDBYMdlS0r+tbR58jNiJSO8mwjX6DapD2mDwpRQV5GAlRF0HZz4xxcXQ/QKAbRn3/tyWLIoEajX
X1L3LBPDSZTsXMUNEDLHp15+Xy1BD47VUPSD4ME/AY/kAtl3odPIrKpJYKGFL0s9Dq4KCEXdWc0E
+NIZeiBNf6nGtSCQIWAriQqpU4/B8OiQT6+VErqSpxJ/sqpOiLnThV9bHGwA0z/A5h0ZBgk5vjJF
7qFA44nLEBcjGlikOxRzhbw31zJZWY02tQKDmMWzgVZwGdyzH0UOWDmya7oW3HViBK4ijpXrZbT5
nSXk5V6bEdHEsTz/utdHGGgGMvzFphJow3h8wc1r/1QiGThsq3ozE9JfuGQ3oavESpauyKq2mEue
op42Mzs7dPGJywZ/eVJD7o9n2jjbfaqyyMPjrhytigiUYG73sJ+vQ03lyLUW90rFAQHGnP/MJbzY
WoN43K0u/bgunOHvcN8kwdHAIWFayogK8TkAWGvZrSBWNEen8D0vR9HFYmC7PJXZtIfHShCOLbft
JCsyZNKPWlqLACoRwcrSDu1CK9vohjGR9L1HCkzbWzie+04/q/sgCH1Q1SQuMKJdEOh2w2rcj7h/
Vw64anS6L3xqPoknqiuNX6+W2E024hmLJgeVTtQgaJ6duvDDIJfYXTmbo+F5SbJVC7nWpOu7EN6J
2m8UCgaYQ4I/e3yVBSP5lK2fkiGZHv0XNZz3FoPuLudTv8MplRcjBTmKSzxcbjQkZ7Vn89IJQ7JW
+zd4U8uvQrrzEgalAtQ/Znfvj1GVRcxaTufAy4qqmB7/t9w/U40o/+dVbj2HxqdCSG/Np/O8qjNb
f5rFxP8cjb3ipU8sMg7CYM4Q2hKXS1ZxG9uGvXSduhz743Z3aMgUgSl7UjOYMAmwfes5BcvbM3ZC
dkv7yDu3+mJn5sp6mrndzYDCmMC+Ly1TtsgYNLXvj9RsdecHPhhwn8VNUyB7AuR7kZUbiX8yln+M
z2RyN78S45ODtQPQD7YDvtlDCbzZzJXwozYkBpnOMWiolcw2o2HNmRx218Bgc6Umv+KiUM6eD4FS
3cWZUfHzO95UIguaqZ5zNtCBmomLaQlWcTZtx6sLl2AI+kPIXfMhMrCbfXCb3icWMX2MQMS3zYxA
xB/MlALXFmecCZeAX7n8hs8mFqRakzFE4s+J7+2+2iUAgrAbVbafqA6s0yB1iUBVhS7WC2mHNqrM
ADQBT86nMI4uwsXa3zrUT4tf2hNL+ard4TMKKPTXSJHJNIwUfX8AiSAU9nVz9zorCJKGRzQehwOh
5Ha53/XQRmacqoxY6OW0M9K46q0nInCCe4QKPL1BH+WAFANnm9Y+N36Md6lPRtFetFMYeU3ukXrz
6jNNRhLrT5uoXy9tgglTw1gLcUwPNFxcnh0VptrFBJFOZTX1uVqF8+RR8CVbeK8YHqksVomETly+
UfzBhJY3DOxeUp5mlZzDKJcCIaZTaYogAvrGUrUuAKlDUxAgIpX8mQfYLP5Ey1lySwCaY1rtpjPa
iFow0Ck4PRLeJ32Okg+WegyyLb8X6KL0yO54UxborHCtNYIVqNylKVZL24EX1PJKlQ7t+ATRuvU5
e2Y4VoWUQsrK+Ic7LqOx2Vt8LYy44spimLD9AMwKtEK4iwabUsOFXwvBL6zkX2b9NwDiephVz7ps
w6JBPM1exPOk3/1uGdSY+5xqKmbz9yjYHGOsppUh+0jchnNPH1MtoS3yJkjsI/OC9cCrUfis5YDU
3xYQ606+ES8tEhorccgUsIEyiSwxLy8nhPaixdw0WXQ0mUPHMl8UmgUCAWG+wUCu5b5iaJ+nYrFz
64hpkxd/VNXd8LIIWIjxcQJvtYqkxid/Prq7deMnCCLNEXa+HPYwbXIB674jFeZAob/7Y3b/oHJF
x5H2eAVl3SB4hP9d/vREi6u8yT3cZCZraaXHcN8bdzcFrZ2DLpp/Zjugn6btuWfv8AE04InZaKse
ohWZzFSmTB74eszgpkey4zZ66/Rh5DCp40p0cBc2grHO41sdGHvYY3fj/lab9rj307PIGpgALyGK
hhIcwMDc1h2JbQjH15YDjpDLJhKKMyPN1HE5NuUjgzlCRlozJYLQaMvwg7V+OBWFS7mY2/QriRU9
6r+5c5JileU/9bVSTsBKjaZsI80JRuy3q3+kX7zBtnUMZKsxlko9sOlQteefCd2qCaFZmLpJX/3G
PT2lpN+5p1O4E3cB9IcEY7sII2btWxHQtR7EKSOK5JY+lQYGLvqxCPO2nToxKBoYgHxadtgEOuOG
VgtMF2br5FIyNcwtM0dC/rZ0Z2KytnvXUdr1Axml40NnByhYy3KbwQfnjclIGYSPNFhibJcMKKb0
hTD8SLkqiGH4n0e/uB3rXsi5z5uzS4o8RiVQoQInYd0VTZGnLPOrcOSKSfYdWpAV9RSX0U/po9IC
NEe0D9cCkF65zKK8Cg/S6DJyhDnABWijNSrDORL7rOLtcPOFrotjbFbALZre+ICgkqIrrS2/2TpM
QOmvuzxhUAaBH8wAF7F4wl2VQ5HuR2s6zJP4xPFA/DPzKdjpJjVY6MGgxpvoO8lQkxrvupc2xD04
fWBXxptj+18Kpko5Mp9ENFyQxG3UDcRBjzNKI28bUIrNwgO+N+3BFnfBGriWYmepEJ3oLBDU0aKS
k69kL7NMSpu51F5fFor+MYJ/0pSBYntHGe8VZ1FR5a6DbLk1p3mqEEyCpCfRdA4wkJzzo8imSrQ7
IyZnbOWvx/l9COYaugKx0a35ck4g+00TXYWRVpupWf3HPBwO5R695c/yy5kxEegegwEroYb/zmoN
PWQ2TRqy3/4n30Lusr/AOpDJC+A5w7UeaoSHafSNNExabjWS5TqAkC+RWAD7q1vSl7j/framiZdp
0aEE1lPBiJc027RZKQkBPfNAuPKQo5XShbsGPs0GeaI+yKzOgh/RbbHFCxkqigAxsFFiaXHrucwf
JV7pIVJul+yeB+yIIh+jlcbLD3iN96Ye7bTf/j9EugO4gKK/o758qjDjG5MOpOULhCnztkEo6yLM
5L7KsCb7VBcGo1gTfZeB8kytOPj12K1LSlonSrw3+iFEVBRXPj50RywpUrbG+mamkwqQFafLRQGz
V/4UQIT3CLIFEOQp+hKm+JCpzlJbcii4QdGfQ4jIiThe6e3esb8MwAex8hpUm5lkIDEqsFxr4cWr
ftLah7qz/vz0tzv0z7uyoEKufUW0Yn6tMLuZyZWFB7hWPT9i18hWTA6Yi1iXkkBnk646PpcKp50R
HCxonZdNfveuCmZpA+8FSpviJx5UV4QfrhZLTTbSViumKVOvRBNzzfH3xUeTSAsIsc0DCJRRPxek
OyxanJ29OwKun+wmrMWxr299HAjwc6gr0P5s7jfUM6mLNNklfgxziWj+1BD95XXytlsNVFjHa1Ka
E8HaXy53TkJA37DKY9Y7kaDCu+fF2UZB+MD7qweYMh2oIuOaQtJkEk15AERwB1PZzu/OSkxEmtKV
2J9zZOjGwRd3piDJr32aOLvQDVOowb9IUFZqCjGdbmUo57nbaihrOiJyKihKEw2CKoJTWtLEkyGz
FVCYdb+Rt6r9zacWF14JwWMnQqVY0xhX4OHfNHzGgAaLJgT96Nawzcn8LecTaxu98hZWu8/LMLcp
v9XpZpMr3X+PIPr4ELpUsaTvTmzQr0VuDL/vxl+PqrqsNsRhGRBpsk3S7o9QgSUOyJes69LnD7oU
mHGZ1jvZaKMJoaYOmJYLbGo8xXOX/muW7CdNhE+QRCIsrhtgzbeMHtdrJJvSxztm7odwupAqeUg7
+odxGoka43Tko87cQR+uzDFnBeCYARLibEWnvubEVqgBYZy42D0x7ZoZ7E5zRkx2bzxuT5ZyQBqH
5DTQZYRv4sZPvf6tWDY8ej/P2Ip+ySWAwfQQk4lEJvmTTFHLtV8hhunGe4/oWAdE4JujQubMu3mD
DZ/7a1F1BF5TWcsJaxn8vRq/xFzrPmtf3xfLdWE6291YZX/bkBoT3SvhdIEBYq9Iti1EpcOk2lfa
E28S28IYIdRD9xYET0IUegOGT5vhdabkE6HGlfePvQzdZDvfetH93U+JEImYThmNdYX9PSSTd8IZ
rpZ1u9AMfRdo2HHy4StdY0LMvlPw9ogBRxumQ2QfSSNEmPfBUyEUc0d8m9I3kPm8qps74dwQ4CVm
LE6LNJ2On2psu4MMlGgyuS+NZW0O2DC+eF9V432Ef37MylK2H0GTkomKtJxysbbFpWVAU5E6JC28
BZ/RbTxZ8vw95qD5VI6uJq91ni5kFXLsnolPlZ531vTRocVurAE0lptHJVBV4CjxfXaY6gV7bEQW
1duzCnJZg/fXkLtXgZ8clBJmZyxFrNnA3xNxla3X2b5M9vrEUPcCTGn/Ixlg5hCjIBB/hzLmOw6L
HqU54tGyd/+G5DtZj4iHEx4e3aYWf7sYOjJy3Azl9g99zz/gFYBvBqv4xQh6vptLNfLtZaZZsnVw
58FBftg08Y+L/3uVvoFXOsuYdwbCNqP23mIZyo/+TeJc5fHdggHH84ZgKKvCUikNptYHVxqgKGiF
y7cxzk2MCxXKj+A0StqxCoIXviVa5uImnFFdOmYZ6gpJYyo/p2/jlnxmNC51Qnm+qJdBsG3YpSzl
hex9KcaU50deb9c+K+S4wtkab4RHFLlZI3tLnVXua3VapHSIYPVmwyOKTJz895KjVJqrfu2+AYeD
cQvWGTXLOXWf8SoNUFNGCOdw+spI/GACuz4/K9gMpjOXQrpW9YB3baXfniA6zdK6A7J/6wxlQ1jk
OQlrg3vMuelwKt8nMqkHDe3oZMjKHKWQNFMf/7DFLsDrw826zRG2wYgtvpztfNymWCoXz1Ukia06
hkpAG0/PMYlE+Fd2ErhvFivrb2Kmz/2Inpa+wWMGtdRrIASZ/MH++nZMnauB0F/ndC0EwtRH4TMQ
GBoXJAkAfV/kLfkmPgaHj6FCAYRnTrLCb/SoaKoFwSS0pbp7y/Iz5uXgYEw7fwp/X/GRGvFyLaUV
8+qiU6ourFxfHUYTk9jx8fzDGB1IGVvUei0A5LaSJWV9AZGdpq4OF47gCmqO1XRWXg9n8/jVR180
M40wl/8P+c0YJUZVzZO3id/LbJPv6aqTdWOZ50s4Ws4M5jF9GQ/QUwpsMW7NTrYEIa8f4T9ojeUR
owH6brKnecmGZ/EQcwY/wepI+fnrm7jxEGI8u9b2mqB3iz2x+RWJOmYXmszMfva3cSjpn275vlL2
JXEwXt9OCCSMwUtYLIozdLsADFCaLH3UQDgDn2Aq0od/zRjy5iC+pXJUAt5Y2LjKU1DasUZadX5X
X01f1WFKJmlvZoE0EtXQpROmu7fdEOcIfWFX8jgiAtipXPalAYFWE5qFsj4MqPUoj1eBTAF7Vyyt
wPGaOOh/opkuyy+2I7/1YiUyU0v+gM9Qu/uAl4NqjHqqoTukzxFiQOCoeCYwpc+mLwnD1Zzk6y/7
1whdOcRBg44q/e1rU2QF5c/PyC6AwSbVDtyBxxWQpsC6vU41cSLF9IDuQm7cscXyLJy5FFnHc8zt
18LXKPlpDNJf4MttdCE1h37huuD5zYhHPXyKdCnrLuTE5Fid3GG5kUmf/bofXHN/H4OFXcA2FJzE
puk+pM+0k1m27k6aIngseGx5DU0uCLlonRB4VadAhP0VKJ1dtGr1QmHEf8k6k5Ujz/DVawOU204P
cuZ6B/7ctF8H5PdonN6EReXfrMO7sYGqCJoutiIGg8IcMm2J43rRBZQIGaorO4zsHRtkzr3jvxaB
Yz443dejtOY5U0L5PlfhdMe6KpRDdPI214Mg3buwnBgq2lgdiTX62ERAgQ70NRW5ovk6lxC8LX3e
aO6pS9liEJ3yFKGhtl+CbIJj5p5v5Jhcu+vU0DLI6/nLvxW7wAOMfCPCM7CMZtqxjvyN4R9ZGKwa
L+1MMyvovYKTUa+ID1CCyIzHDcAU/voCHFdlW+GND0GQRnvtNPzmP1epYuNHeabNzqHs/7Va0enC
Ik3RXZVs1WbpEtlkBORdBOn/lBE/+fzgx4qlt8TOPEb6TuVfcs9oATPC1OCK96yLf2DN5fv7BlGM
6OUACNMjpDF5PMamlsZc31cA8igyG3DW1PLpGv2rZ5Xm1D4hFPXSupM+ku2XUvzneEVoZhQjjssM
eqlFEVQYAg7vXEelJYFlNNi44GFBwOjtPVyIiHSHZ/rjqEFGOyCApV23d0SZjq7OZ2SZw9hQas8v
Qw1XnXvhiHA1TvZm4aw5gKBTTjPfpqW3yEP14g==
`protect end_protected
