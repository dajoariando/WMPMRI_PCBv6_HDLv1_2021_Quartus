-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
HDuGGOwnVjUva3PbBncT7mzl1rYcQGt1MWvP58tmdZhQaKaDwbdAv5tlyVbYtrV1GHri+uT9im4z
QMmWSQFEdxZq3f8efBRq1w/xmvaMoPhBi4z5HQe8X95kAWo5U0OdAxp2hFckjhcGBwuWz899YkUE
lfbI1MEgXZijeEgFU9nP9Bz179AzXSpHjAAN05gJ+zOuIqbGI87zGNg6gPYLWyXomNchs5y1IlQG
fQG+t5qYKd7GHFyG7lIOsgt7S9GFdREVN46dKzN10/rdoRrqugxsOKr0KZM4SVQEsqwhDHzYQuee
q2eI3d9mA2qJn/+3XyOTsQMRhQdw4MzXPGd7YQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9712)
`protect data_block
XhTYuFZRGyvFuG1NVOGCN6kCMIPhfrCDMGzMd6QY6YHESiEvM+14hjjpf1A8kjHgk8tEEVct9TjM
sy/V0/ju7KyIV64G538MIaaFdim35a6sA1nt6PdpmuUUwXL1Y8GXmkbh5B0aAoIirmoBM40qP8pD
fqDoaVC8+hN6qqUe7M8juQw6cDs608Ve0Kp5lKMqUjwF57u5gNQJwwrU0krLqbV1VQi63KGzYXRf
8iBVFZ82PhJGMdoHfO2nhZp2DJS5hmRVKaxNhj3CRt48+ag0S7JpNiwDmLhrPHjyXJuQMIexB49O
P2GDvxkGwgoRk2ClWbsZMML4Bv1JJINxFWg1EgRUz+d8S/diFMS8YVnyOjl/t9CLQ1KXAvg6rbRX
aua1P8HTzu3gHz6fc28Hvvjgojw886PoyfX0Uh+Ep/33X359tp8bL/NsQnHKqExdLT4g1rA25Jpz
uJb4smPi/rX2prwDzvvTg9e6tMyJKs6T8hKpXkvX7GywRR51nQmKLlxkfItk4TZ8ygKOa2yZskxv
X9sph4bMbdIczJpGlSFWtxkeeHmIh1iSF5XqG1o53D/GzOeYKNNHoYJU789htuhUM8N02yN4FbuI
f9nEoD6u/6vjMlvGIGlWNf4mepI1aEixUPa8F8eUeuiVz2fsV5eqznz5V6GbzPRjJ81bMfJ0dI2n
Pr5vp5UYw9jRxgqSNaaONXmx098yPcQ5GuQ2uqbuflUl+4CI8N/hvfWfMS9/ZRY6uffIZ7Ab9pQU
cFrQw851qkZfZ4tf/HKtiD5iVbiiGN7IGmjxtIlQ2Iyi+2O52wuu4UlkKM/syvEDQ8cukRJSCAo5
t7Mm2DTPLwo467ab3LhRUWxnx3wk+Vu6zhnxPhIDLhMt6rcJorvAvHfnCdys49gxtqHZIQOJf4Xz
FYDBcyY9aLD9yqqci44TCYaKb8NvNvo45nZGXpXSwtZCqaL66B+VPkcJ3HrsInXMNo/+ShPr/I5A
88AsESrgT+2/wzZKbOH1fgaOTWiiSan5+BOCANImp+DWMnar9wvzc0WloyIY+MnSQpNrBKvRMjIW
TXmK7K+ZjEJP7UVQcZvzEsJE9mTVyCsfhCyyBjN+REn01N10ccW0opbcT+FoZ5fsva3WKNvq7yw4
B7J/A1yu/cfBGrNPp3Kkfm/A6f9YczdAOnRWxQwHaqy8WL1CJ5KD6D2yR9HvVmRKGFAZbpuQ89VA
zqviYS9VT17WWW9Yl7fJgCfA37gKp23COuymCckxkX1tu4c6bUii04OggwDfNf4829CyrGjpJZKR
Q8boO0EQqHsGvQsA4nCZdi40mJpejtjQHLf+Y86l5GqyOkN/t1X5yLQYZPKamHRUMg2fB11Fqk7D
YOkxGSSh0ADq1Cbd6RAul0rMJOpHRcf4qb0tCO5N2JHGAeY+sqMsETCOQ79kOKkswCltozXw+fmN
jLmmcyg8Tpx1bGIg3/nDPk5P8A/6ktvX6XLtZ77jRlctc/cOo+STHny2yLniWQMoXRY1LSr0Bhkz
A0A60hG9ohyZC21MoxtCtL57a80e0srigHFHdjdmmhPPBSiJNPaFpiCi25PrKrHlSbZkaUAWanRU
7m6IgPOw7OlIY7cZ/4CNe+4SSs4sM0JFZher0hLtcfTaoGGUVfgtZfqqYQcG1JiWBhNvIsQaFZXq
2FkFekxpe/28Z7q+6yvBlTRlvbHLlFMvebnpJ2OCSyvnPCp36ucjFOIluLlq+biUcwd6cdf6S8IG
Ly5QUFdMNY/VbmDwEJvbbdNuABO94IHld6X8u51z/6apEm36io+8rLhFQMjeojCWpaw/BGmc1Fus
Qkqsr/TcvEkHTEE9PjA9aeViQYxCSfo5lDPdXjFVWT7PsK1g5ABcey2v87GWoSOMmMeXCX/HPbli
KrwyWNM4TNJNt2ZrjipQQAovVpzo/ZpW0twuXdpB1QoxhWf1zGxXdUdhdTPRD/0+3VB9sOaVO8bJ
9y1tgTgzbcfAWNz5HE7Rfy3RMhVHLrrAVXBz5M9iNFjOaD9AR/yrxWxCL6rWp6igCDEzzuNF2xLN
yr2zDmWHLKo0vyER8K5KAm2aIYzXcpCqX7ITvZgITRb1KfB38o/aovp5YBK7vKoDyaCYd7emAIoV
TktYzlNEncgCbqSBgj2yWjNDgoFsTRU3Qd5v1DQSB7RTxcpZ62B5WxjQHmwk2faQxFzbTo9vpm3s
Gk13Zr7OmV0CUbu9qqkc/CrR/9UTN48DweiSmkoWnfA7kZkCxM2cAjIm4ZQJjZBvRtpbjV/X7jBH
Z25COStyKDU0Yaukitn8wfuUiS56rvx4Au/wlfmQyp89A2YiVmNXLwfmt8wjdQtPMjf2cT3r4tRE
fXHBB0mhvu5jUEjGFTa9+vjUFo2BjYmZ8qfmYha2BKHXcz/eEgbGRR7+dWBuwYWNx6wvXg7X5xxO
2eWHhQ45Szheg0O0Hc2douDwazgGM9dNc2+jhNl0SURp45bwvY+5wYHCZkSRt6UUdRQ+K1vugwud
2W7uGh4gKfmrM5ZpFsgia6WhhXLYi8p0PW2SSwxLJrJaFqigWUusQbg8yHx0DyOAMSUB03stSnVG
kkMokt1dybQ3gUPvnIl/NuzxzjVYFiD3cI1ktyEF9piJPNgfASr64bnQXzqYnRNNe2/RjhMVm3Py
IgqZBzNEcU+Kz23ujWIrmJYooVocy5LHU3KZNNaKXv/5fEqrEz2h8Cpq08v7o4pk+c5zGZ92wyGL
Hff5qlK8yJcJIiGxvAsoEf/r7ONVv+O/dz0t6G3uVjfdAXjm+2XWEwFvYBgrrjOQP2Air5SN4umW
BIfBInqj/BE4o38sf2zoXau+LoNYTC3AA4+PZnwJIXRU1zBCX62NJKBodQ/BYTMzTWXMPPh2dy5v
Hl+e5WNA0FF5XXbQwdDssPOJRnqMZHUJEuQ+jHMmifVEGJ08QMhPhZfXXgA0KdDOgKRiTUFnrB2g
S29/iallQHJjd41LQ8uc2GTmWwSBNRn6V2Qj7ZWWSfVDxANh10WN5cHc9oENbonvvoRToxOcEKHP
vrggx6mg8rf2X6eI24nsQNS4OhTz4Y8lQ6MiBbQdnEAreo7AfBplh7b4Qs+zTHMWfGEPId7970Jx
3fSPYEijmwGXFvj6c8fONXY/Khz2E72LX67eTyfyj8V3EF6oQ8p/QS/YDrdsVoo25EN+jepQgAeJ
puWGPUESsqioUJlKkAepLJeIioGOpLIo/ezdyJnGMEWpdQL/6xS44h4egz37L3fqjW1C8hybsP12
L00BF6Y1c7C+rj6FarZ4B9URwPuZlaSnWicowQuXfTmkjnEtQqZaiID6PrRyTauBTNn69sdFIobn
xC4cDxdJh1g2Lh97o/WByTIsdcr0yue+eP36bLnQus7WQqSQp+nLvi5XJ4tBVt1WhzwWvN3xspzi
T2Oy+t4sgOu+KvtAc8kqF9Crd+YAXZ18QN6f8ryM274JBN37JBfY97UJdDvvp5DLqyrQtk/Jjnsn
LGIcA3Qpx1pr5H6erFDiNpGSF7eCy0rDzxDX8HxSpxGBGR5ds0knQ2+qz+BGi7D/O+R/3Wy0yBBh
NP+NCyD5WHm0+ydrRYxYjoK88ZZT47STahlO98g3MEwF3jVNowXQcoca6cw8HjIXYFa+HH0Z+uu3
3bN9aJdsbAL3ak2VZoVAWycdOWxWeDd5HHzfUgea5JpTNDBIoOk1Xph7eYZQ0waW/Cep74A7Zj8x
GDfp846dDg/qipmDgGBoGqAtpb6Qb09B6oHvShRhuuHLbYsV7cPEuef7pBKaB3wCnxE+JXFL5GXs
+pqBg8QOUMHo/keZ2G7M9CflfJ9xxuwr/Mt1Kx3qUG6IY066jKpEdvPfpcLEbo/jo78ksCvDi1A4
u5TGk9CIvE4JBMH9ZLs6tp5X4kpcUPa6SPwmNCt2KAluIkolyxqvDSXowIp9t9cxP74Krx4WSim2
AeBGjqOYEX4Z4826VWs7IdNfn/HlBy6AaF0t61MrKITPNLNY9lnmPfu7tdulXrSJOsVnxb6nJEe+
L88ujtGaJ7E2cqFlNByJFKU3ftun6FexQ/ODpnuXaLZFBm7iI6QHbX/15c1b4lYGpnTpO7UHIG0b
Pmk1iLZ3qJJ09AvMuS80R/VnyFxO8hBBDZu2I7vlGFoh85T9RvAxO7u2fzv9+k/vFe5j/BtWpIzT
Y3Z2hQ0A2/2ijBStEDKHJT8P2MbS89Oxmbz2111kFeH/Oc521eKooAqZdXDDsJoEKh96/l5ggrry
WvTtaDlbLgmM/EcZ8EFu4NNsXjSDYmWfqGd/Q7d/Ev5tDPO/DXOaMLHrJExeQx30dCCsIyaBlE/+
maOLnG8gNW9kls/5iqgt4X2ccVPZhaf8HQ9stFYTCdSDucmb6lGdcmyJ04lm6jsIUOXX+bkQ2s9V
Qudhl5tHWDYiKsmDwkb4GTnW+KD41sIhMQkOn6OAXZB/R5pJXi8GSbr7u8qLNW4QeNAMADYYofGy
QgLK1oubaOY+1PLABpWHq9h3paVrRLaAKq6FB4fL5pp9rWbcgbfg9SUZl81QJUnJRXVpYHToH/In
NSEcXGjbe5mQIoUeXEbm3sy1rENJKAv6qB65D9f6N/UMD98fCe/rcWXzFhTGL94Oj2cfvMdFVSgf
RP0f6kggNvDAiAY1dof99KDezDiPsGbGYXjuaCgEixLyilJ42USIxROF2SEwbS01tekpf05zybtp
M41AFMcLlH10v+kpUq7qup/BQ/1uCD5Ql8LF3pMGKk3aPrggxR82Npwk1C+g7Hcox9fdtQgtxa7L
4k0Pdgea2We9tM6hgAjmALcoYEEz2JV4m0EPT94quwYxXe1uGzE+ihXNZ3pQsN+ZOMEmt4KRR4IR
9ROrcaGkf42nlHUM/AvrfOdNR0JZ6nBV/NYA7P72nc6JPSyyfO5gTOSxS/CRkauST+rebWxbf2R6
9x5J8h1DtA46huA10ux/ZNARD17W5Nt08I+i9eHS5rleHDSY7Zy9YGFV5sdC9P6iGKRRfL0INNyq
m8/bhP2embWNVD5RbGk4bcKeUNvl5CU07WZ3RUA0ZAqaPJFm1UhwTK6SAz6O+v8V/OMSJvP00Q63
IekNZrfIhI174DNZyiwr+wTAbNjejf3FWpx9dQADVocYZ4EcIPKL/H7esVb4xbALbrjGjK9GwU0H
/nAI9bAOJWyZ7vdz8Blu6lpeSPe7z8YNZkThO98atgc902x4Nw6cwMcjmaWtpNgm3k12uLIFPbuv
WfVovWKiloOV5G+STsdLXQaayf+1VkP9vag3SXFheHgWql5/BMQIKkaxgO+nKbhmOgHeh99Idphm
bzGd6np5TIG79gZVe1Rf6E2wDYhnHkqytUJjc3hPt+gjQeCom6FWQ8yebTFie0L9aYo9rbZW5SFd
bFTSlHZC1i4cd5ch6XjqIItDKT2FJaiNEr0pobPA1Y4yVMIqJOeGUcVtE71eCNz93++HJk4LycDE
V/YBONrZGHA/OcEpq4PZwjB8roQ/ZUflqFhJABJNRRMytS1t+54K5qNHxOnJt4oYGQA+ud34aWBu
2gWnq0qfWsXFVR14CeOmKt0E9ZzZuV78sDXjz+hBoHx1E5MzJn4Z3aykiD4rLQaPw6VemxjK39xT
m9kBjyYVRLsceN9Cu8ZYBpjgVzBOKziC1QrVh0KEvxsqz5n488UyftTqklmYk9uhSfZmbqqM5fGH
L7mEQKIO/IJTBGa7HaB6ti0DgV5Nvn4Q7ZZP4VziX6XAAcpU508SC2z/HUqQkYqg3R0Z028M9ztO
ijkBrF2l9WAY2OWB6iDqw5CAei+oQI92vIqgur6WHFthWY1eUdu/NNVs1HgSgGQBXz5boDWB8mh9
1Nh11jv8UOFUqW6STc9eMzgvlXbgAhBieJPV1ylBD2htQVdSBErrfs3bPprMymz4MyU5y0rhkZv6
mURvDksYOCCPzfcZpGrH41qrh+ahQSXiMrZT1/G+97chvjLkbXZtvJ6llKmobljCtXQ87J4gOaye
aQeoJ7J23yL9Mx+eQrKSkETASh4Wpvbb28a7sthu5Tg6boy02tvqC5KnYKycSSkGZXjbpTBbkFTC
r2GxBEaEjA1g1eMbKAO2AZYmfDUO0SdbreTaGLUm/gCEc2EJ4k1dEgdPAjHPY8iLO8N/Kpl+LsOK
4VObrX8iUIDcDLrUuOgQ7oEjqQgWt2ECO7dDe3A9mWCJUIkK6QR2J7X19zt3N1++QbqgF0Fl7KqX
d1Vwh+KE/Ygz00NibmmHZ2vrwq7+xPUNQlyP56n4puJSB/9sDSLT2XXo1nTIw7JhMnHkLOISDDCN
FGPLDojiM6xTYeypZ62repdzI4oPk10pjeNPJKJNkiuOZsAz6p9RoXy3ba7exCvt3gPLBaSLMDDc
1PpRPKCXGW6nSFfIRBERh8Vd29YYhlC9B2uVfCxt8kIrOaZSSAjZ2pdTjvzdUfX6a0cFN+UAKfuk
fDNdvOtzbYY+CHujZqeG98Zk7+4XnA4LX6pTrOj8OD2w0AIaicpMKPy3HJBBqitL5Vaa9o8A6FwF
9FjdlLc8ccuJW2H7gYAZsbm7RJ0gIFlmmgmJkNFMxkOYwyHPlyDfhVWk9OlBxabkbxJezdIBauyl
S9GqfLXEQDZ/TGKNJ1OQGYS5CRyq90siEgg9KkkiDpaWyS4gctvJ8rHNWB5C0Yp1ZNr3209OZlqD
WwtpDebKm/NregfrCtgFOJzKdYZRRjIVPAeYnAo02GMvEvtfAogiKU2Z1L879IL3m88ZRf4hTSuC
Oj97w1641oCDv8YiUVhZvInAmuoMDZij9i1FexfkUIG7s7Ao0+BFhDOJKfxDvL0cj3ryXt0o7+RY
/Gtivc1cNomk7Y8epx1pzGgS4cmXS/BBKk8Uvk2kkJSdWCtF9zJsSo/tH2ZRnbHIEKadNgvb6v+D
AOaWCHHbuq7jH4EdqO8I8aQ3p2ZCLjvO6/+1W7HUJI3YgREqxOlVvOtMYYdKr3Yc1iSK5cMhzIFn
CrVBhrrPkuIst8I/meOeyS4GNGRx4ceOQtzmW2yd6DcP1cB96GrAH920NrHTMVKPu5txwj5NO8oR
S5i/OKn72h4U//QkI93YPKGs7dSCJMlSorB/0zcsf9otzH6g6WmQFaHhhp7jQnu8IOkd2hDWYz4Y
uD9GhIcvGvpLZbLeUvtVSfl+iC1nE4b0yc/84HDIAduWjte82leNDM+00a8Mi3u/tFjYbnAH3xDy
8Jm3phhArDbLLGKNBVF9Clz+kLw2idp/HPKKn1QEv37NUHilBQpXAndElsejzr0q93HTn6WCF4Zy
Ao3L//Ar4T4Ps9QmDQ6x52/K9U5PQzjfRAMtCnoO7CoO8XER7BJ2G8wd6Zedrtj1q4kFUeIwOXqW
LpsikLjR+rpdmJvNzDnypJS+qO/uZDWWrocgIoMtbnXWxO72H5qXvMo2TW2Z4Rjzanuj4BkCUdDS
Vo6daar//8+9exBoYV/pRTZ0wbGMoQmrtYfHk50WguyAu3Nc9feLJCG7wpVYOwbJnIn1dVpIOR9T
lkdFRYoBSVaCnmigTJe1Iq+HOK7TUeiyYt3xMr1UXj0IPuUQOQJnUiio1gVlF0HTv+KsMBtnUlNG
6C4nLVk0eo0ypxNvhQLWdy/o3aYA5B+P7be5Bmb3fj8SDCAV3urJFQKkS1n1SD0LRc8B6/eBZcmp
YxDQJWg8+W5KtTg+oNJv+gSqwk7Hlj8u2kSHiMMmEM9V4oIyiFt+J2a7wX7+Qb0IV94bf4mxcLbi
VxPuw7zz3PvciNx97WBpfzskFAUH+BqybRI6Ep8WntFA/nwP1h6pT40mYuH5cShuWkcH2wTAQHjC
2boaItwWDe7vXdzcXn5zsJSnNW0BJ9ia5FbTHCo64lqXw2P8cb4mCrpmySFwPr0kfv9pY81MqAIC
Bi11mzgG9y/nBbxvcdjzRHumBfw+Rd9rRwypw1L5SrfXUtRCbZ1rGk/LOml/CHOTsF0kxf1pCp81
Tef4sXHLG7JVIGu8LXqX7Qw0Ol5d2tmfD/QI3z56O2SCl9naFQnfowLjGrwhZOZvk8QrIVz8/Akz
z8m3DUBej/8FjAHpjnN2GSUdVcnUtSs+MJ27FWCJIPXU5nBehwCHG0e/eszd41meC3JFSFWNkr00
tqDl8mnjm94t+TKjI9TpFY0z8sYxwl2UCspzecjjp1PF1Xg8U4OD5EYPMFHN4bXgySDFgQGdS+Tv
dHfT5LOj2zLW/JJFsHmc1lQnrVZQX0emLMef1rDZe/CNv6oi39WAe/1SIHkXHMMQc2CJcvdWDk3x
mQv/4caSfGxzLhCBNUpklga8uBHwXIbtE3y5Tswrg8GP2WNlXxgLXt7LKYZnyeIF6Bl/LamAgq4z
uj5D4/apokT6Fb6rLCctz2nzKHcSvFsQIw7xMFWA9x72SOxmlf4OCAF+F4Caa3RKi3LHzqg15HKj
cwbfw9vjpLVTGcZVmBSDc2SHmhd3rjEpQOmwIKcUMeMiKbdDscU2l5hPCqUnKFgCnaiYjxgtamDf
vfcXaNu5tny4uCPsq8NUGH8z2ReyUQXfeiYnAcdAqwcgAyPyyzr5bP5BCRTTFwXTnAlEsRDxUEfG
JpP548lSFejG6U44pTLnKAfAgyOVtTKbFPieixE2K5/HmXTgTSYQ8jTv/b9VkD0Tf7nwae3daSYT
F7LZLP/LMZuTb3u4tPWEFtgstlrEj/Fa1TcZ3aDKlseJkmNxxEMWduRyzRysXO93m3ftikDHYWeb
GmJUy7JkUW6dAixikJqlbxZgoYJCT2uxhKeN7mIovn9O6bH2TroKkueVECndQFvKAn4Ht0ESpAZU
i154WJsyJ6MuUgmToz38HVNLFHGFUE63iIQn4ifWTb/+TFJGEjF3FK7XMJeY7EQEhkSSySUCTo6R
BojOBF27/5uv+LsUnIGMcqrPO0AKAWFNSDe7cEw1iBKfEF0l5lDDNzEs40Sh7z8350FyTwjKqnFz
/9J+C10VfKhbqCQt+cJwb1+uv965HF877tVyiIas1tQmXMW08lCFqIdPjqpMM8u8QdaiNG9oeRse
OpLj9PZmfdbGTxivDd0dB8CIHSeIuFPXnXG0LL03yR0+a3ibhDETcM4/m7c1XP+y5biZDh/55D/i
G+3u6dcVhpQxqVZwO3qr2qbYbVtRtvq/NqRhxV+3Ci6VYVN1jzmZHbTTKqCna7RYsFBRdeSljijP
p1bZ9uG1nuK/r+Yow8qSy+V/22d6SgSgKHpu5gS8i2IdECeXuRTpgfK8VZAzjtKGFxM1AHPk+I6/
97LKSQGfrfpogD+1QEmKdKep7ygmt6r9i/zI/oN+84oIrBdEMC3d79LNGYagU+nUbk49W+ZNC/aF
RiCfLBvugEz6i1JjU8hiAjrD58rxmkKn40iAgF1FQOhBGZd2Ti5y+SS5dZtqISsOLvyZJlt1yspa
QIIIA1HbZGFX/4ZBy4ZErL91q+KYpx4MopBClHy4YpITYXPWzzcPuvpdvfH0gCVhtzAAc9jkVdKz
E8RYZYVwyRFA480bI7yIq1FTUDQYs7JGIxXcXdvSky1z9XUauqY9CqKsaheeHp+TtBCIxkIH6tac
3QdojwtMBfh1KigiS9J53FNNErK5iqJtJwWRIyBytZZB9y4//rZ1LU4wn2GyPBnhhIW5C1VfGnu/
5xSutebloy2FumQVcqxu9gzBquTcYBTgyzgjbsBkgpNEMWbVAUdBvSe1PIg6NXld0wUlY6jp04lB
9FMNMTR5YVYRdNmRyBSBf0lckFyT87OvFDLsDsqOWYtsGiGpCutRNqStYjZ0VVaHB+Qq05w4NzcZ
Dt3a8ytH7vCO1D7TIs/7dedG82ZIwp7E6NFott7vcS41vHZvQkcPVbJrqSzWulRGRlQww410XTQH
hnARvwzrYXAkUHTeLNw9YWwvGjdZ9nJG4SE4qIlpZ5fwzUodoZ9lXxYYbOXB3hs3uNDOKdp4UADg
LUiJwkQRe0H2/zOGRSL5FeMrl5PzXHkAs6yx0bezloLgnByjDBLhcnSY2OV5ddMZNG0xj5UWlV10
MuQfisa4DfMLf2AmFpaUQ6TxsdXcvEXysx1Ssh0KYVs4B9JN5v2OAPfSnSJe7S5U2K2aHrFDPxUU
y2rCVj881SVqVkImnM04e9R+AHjAWdT0WxqVdhtChxHdFQodfszGz0F6Luaq7oi1IyGOBRQ7moqj
0xQ2+MFk4upmsQzp00fiXkmNd1uVtXWjRCRqTmgvjYJEj4BIO3Bndwx0kAxWWOUWEzmbdpN+8nSL
7cZKKVEgUbbmnjqrPZeDe+Q0VFlQEM5Nqk4dStliToPWZ2/COcE7QSAQP8gqWmBPRPNZFhZF2chb
SvRPCzgbdvCKwu7bKEJ8m1MJ3cnnEO2eiILKJjZEfX+M7l5jGoN4vSWPnP4iTzleiClF8G7lr73l
L3C/S+tlH/2hk6eEuqxpJngG88KSxIccaMP3ptjQKLs7zd8aU+kcRbJoHBo7V/NcR9sN8tciB8jG
KL06dO8unjJLW+jR8KPEyrVPN3ywn5BFbwYyToZ7b0yLwciFMY9eft2Z2Pr7D41YixCBZ/tRPBt3
go+Qb/dcBjtSzccdaSBJjg8puNXSW2xoQoKgo/3HJv8rl9jWJYSFFM2PEP4GIjGcB2UjT4PHB4bM
g/Qqsuw3SIGdxC5hQTRbq0jOmndzsa4ASqCblR0ASPeZoc/BURpvqB7y4b8bdB0jr63CzNVuqs4i
qhwblIJnW8kxoGMaql3kerB3BkEUoY/PSthNlUI1RejRDcxBAOqL3v4BKLv8m5Q40pNAKwgex4rv
0sjF5VxamvWyNOOZe/Wxp/CO4n4gH/ceJPnNrnTvGn/lNnPtywJwFtEDy+VnuGb6ub598HbTZo6t
FHgde6eowJwEf15AyVIZ/mXZQ7tAq/P9t1a/g1dV8vjW1UKt7EEegc+0Pxk6BlBuHxA7nE0Sb9HC
w0/YpwsaHldzveQwer2IncKSy3ietibJJozgD3RyRTiMrAaUYBBv2LU2UBA5hUyDOB1DpMSdBslk
I2PasI0pQzajibZr8uCGl3EjR//ojbMf9qllcsQ/6ep2PDCkQOCQYtYjCYz04Nxq8bmTuOG7qHR7
uBBFL9y4RmCFkweRRQnq20cNn1v6ZknCpsB+XtKvBRAGE3fEdVzq+BkUMYKgruMeSbI6JhHX+gGB
gQjo+P303E1jhBg0FJUHZf2hNY16IwDCqm9w0nbprsuaEFLTi1Dau9H7Au9Kq7ZYPwn7QX6RYYv2
DqOXAx1I9fF0wCHa+Ps1qaNovbXNizEshQZTrFmz4gxCiaopt0K5j57yIUpZa+uJx9UkcVfQZYOB
M0lQbKL91ui/eUkln44qwmO9T7qvqlMnRuTM+LwPdG4kf4Gk5c6rE3MW9hJjMs0GAGFa60Id/hzq
YjAbEazb4SVAITNxx44BvxH9jt/8xp1lFujcoCKG0vG0HEWY1kbhNA57PnxH98CgWUpnNigEzzBA
Ov0RV4jgdipU2Km4xEjiLrG+HdgSzKwac4eBG/n6FM9KjSFvwc54wOVCPRGRnTcMB9J4MYBNzzoO
48ok4Ed3xlU6hT0EDNuVYJUa3cJCU4mgZZ4V56SlKG+emn3zbXqG0/TZApVVf278czHtMGapVF7g
k2snv4KYPoE6nmLzsIvgQSarR4zsNubdBR4IDRSLpOm4PedP/PWf+7CYzamktWsmy/YVGuzTk7ET
T0KcQAinSMt9d5ccB97jFDtt5xbWaBamI2ZFbieAUIF1ae4Shvmg2ytfljP94belNttX5EY4cNjk
RjkIV/ZETyABoFX0E7ApP0Vhpi0G0UzwvciglrXMQnwbFEwIn1N9jWwQ+s1ELTp/pMe35qVCYEfS
b0Ra1bf7P3ngAmI67JWkk1DAqfZLhnJda+QJg4KJnTEdBZ3G6rLrKXzwpNrwyRfkxhNkEWJBhvHN
gIdkzbwxHJ1ZMdV+y7VgebS+iygBAV7Tsh7uNTo0WI8M8F8mbqEfcCimCfYE3gFJN/6rg5k74rb1
CLWxhKk+7FkZfPnXPc5qvER/hjDCge7otso9MUp3F9f+RY/ZV75dzv/Q29M/D2hJ+qz75986cs20
wc6D/yaAOh1vpmfCPJNpPjblKVDaNZOjW9aiWYEIUl7edg3jDw4iIbrr8vK5rW7PZ8DfGAkymTnd
wErAOm5u6BYRYO+s/cpB1U/V2K7kXp2cytTl6PC/ZxsqlQSFp1oXsGdIvNl44BaPvrxTfixeLFwL
TrmX1gqfnIvMJYKlVvxb8VN+ZxRrK06K7k/0mpgoc+ZfyTF/poqBOH6k0tBAR2CB6eAPV/olf5Jl
vo6iQVTJBtAqR4QlpUdtu1RfqgvvI+ms9exXkmRE7fQim7Attb2IVVavR7fmu8i34mVLj5zojNtL
Et6NqkaLpnpJ53AKdjYz6jt2C+tner7bQzHN/0wFy0hM1kpf8tXqwxOcPALrwiIis2oArLpSoKAg
ti+iUQOIWbx2t53q4nMnSH7xfRvO2Ys1vfku0hx12sDdoL1Hcr6tSFmGcTsQcAi9mB6KKfwtjC84
K/9zGEbAs+Sw8Z+7KULdaAke9ugtloWzIy0jsjy8CuD7xxkQQ4+93EqHeq8QZIjuffiuSYkRFoVT
YSuCo6T6qb7sKRK5+3Km8qzosb7jsVFwsodpFdIZqpqRluwroxFWNDZxhVIlaiET1LXij8Y3ztWy
yGW9CaGdemqCscBg+seAtLd3zjPbYxGBDtyJEUi/gxpqCsaGVSxwVxkYQU/Kb5QFJ1Lc8iZcZDsb
PymNyrNT5K0cPEraiKfgTf3i52ejAIQqUeXCFoEcaI1LDEmZ3VZaGXLh3OARswI5GVdXDI9ztwQT
EM3kk3lx8Atc/w/mgi5n9xZdKUEa840dzPCiIw8MeQOxkMXZbk3GUz+bwV7A1wU6dyOgUQT5Z7pi
5kNVQ2Aw9CVcs1lKvJ8EEz1BEpQbNw==
`protect end_protected
