-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
bQZUHqTdDgJH+Iuma/nfBpdOOnP8YZ9Hds4U1cTL0GTME+MpFqAXuKu8D2stmKBsOnJ2BxNd2isC
TI8FdrjRBWuQ2Fk085vJgCmZXKGTDhNOc0owv8FBqxuX+9B3RPcLMxX7RduSNMZUhI70WKsdKHMi
icVz/rFN/eGsF5wgCkve9rSByr+0MwuuuegNE70VARtpZQeJ99VTMDrMNzCkfPxChNAupMg3SMdP
kzeCiomT4MshaKVOqPtLQ1VpNgS9tvbp0DTHKpBIcPQ0ltmhmdFAwEyem1DRtVtPoe7bEsQuote0
5bNDLBNG1b44vlBmzbyt6bJ5X2x1ljJqKD1vCA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 114272)
`protect data_block
lV7BWQLNPCEl5GXA97KUlcIjd+AIDqhggGJxw6hi6a5u+CFP8VugBnZ0tmUxdn7QnLKUZDM+Hz6f
olOjzavOTBZKLA7/3NcMXf4NBtoRDzPCaBf3Hhp5D5CZotu203cy1y3Psdf0A7q7QKxMHJyAgZI8
fJHtacd1xXZ5dMqYXZOtRu+XkBRR/aicRZqRntc7c9E0Wbhl5/lB74QE+UkhoQaEjzWjR4LkxN4w
cgOlFAvZgQqa9U17s43vxl1fdCFqjWDCP70B1TIRn4aBBg2e/Ktm9sRcGA7L3unCxGRH/ffDgsbw
DzIWpPjckFYTFjkLIKgl9gLmUIrAK46B4wajb90UthGJPbdYQhdzZhmCH1trhXoJdBdGcFDDPgPw
Juida/si9PZEII+JWZ/YwC1x1XMEM0PwGM/vjpASJhAYpVKJkvnTZDEt6h/i2YGU7V606ErF4LEa
pWKQGqlqwuSnbiP8fodJPxrloVMRQc01EoEe4aypZl7CJqLAQiwQERH4G2Fc0Ddi1w5YHzdCG5a4
1P6U+dvxYTM6FdS8xpViKdZ+nstVsib1hnm6RvwwagdLIHUuUgHNQf0yV/VCC2VD+PLk8xm9Dddr
OMW8S08tSngTz1/Cr8sPNaoFFaTXs9D7ytspRLMX5ACGziuDpvqrcahdw4+fRda4oL1LC6Xf/WC/
vUYU+kXHN7/O7zuM1FzrrlTH9QG9oZlsCl198v4bI9qP1JvX3b/sSUbVWs1evHftO9q7p0F2Le0Q
2pB6/9CSGFpIM0+CKEzsmAbTBnrGDpmF30mNSFJQcYIEI5/GWPU09qhcUC8LlPxdGte0+zVf78/f
TsodSljL6mHExvOBMKERuuhiJ7mr7ryk1de3oKoVKnuGBp8ml6S6x5snAw0XtodIeiq7BvIE7VWx
w39cWt/ViGGu/8sT1Ks3237ey8xEvh9Y64QOb2/SWRp5Y7pc6EqXePZ+mMPsHFehuwEoc1im3lc1
D+uGV9xa7b2wDV+HcjHgP2+hN7V+cI3qsk2o3GpPRfrWkeKwLWESJzya+Sffy5XMVMEDaP6x004a
uNTtIOG6Hkt7YeQFdRMZJsFge3yow0GVuqtE2zilPvAgrFyAs4HXIfgH9ONBl4HmI7ywVfyXzlZb
YVj5tTeYBKUMIFAtP25OXDqfmTAkpXHQg4PGIFqxQteGVR39SfWxOIQe6OJ3Oa71/F3cMOW4F9Ol
mcEZ/cb+7WAZvF7dpMr/vguosAGZYId/ERJ49MDO8YtuP8xt9slrFBeeRR3uA9zvNZru6Iwael8X
rDk34A8J4B3rdVq1e2AQbqf59EO+Lnootwn0gFFAilutd7Rke9uoO3UNvbRVEVBza6Idwyg+fkvn
fwMltC4H/hPEu5wz0dGKZZQtTLwQwlQn5gr9uWUiWvId9hm2/jILGWDXqSFipN8xrMM+Ixg15W/A
46rw5exd15SULjkdtnOFjW84QQX91WFYSgGN+lBcsBB7SvqdEAji5bJw+78tVbaZoLMPgL8QBhAj
lwD2adMHy8d7v78fw/Y3xUrL2t49SXScaE08d0hXeUke+lyS9p9itmfgFx849D3KlxMz+RAsu6GW
gbq2p5fHdaVx309+ipjt4vD4qZH4x06hDiXYbbT9YrsYYUdjfy83ADPi4HBVDCntYiYhu+O/CAPa
bGQpnB0DoBC18iKghQJAGkAPl6OKD8Nkf9qY4RfoxUlkBetNvIDXpl15z3qw2V4kxFljHueggKij
jDrdqS2Bs/BClL/VuCazmMudkmlWo7fa4ZoTkmf9565ebPJ+4e9q1l4CJv3EKOiwfFFhEAcEM/6S
pxylfzFQfRo5c+a8kDZELtZER/b7SHnKLFv2Sgy3yBxEFrrsGhG6eO/BDk8eHMImOAxu5HDcgRPL
By0glCuqP3nB0WPnFxpKSaz0e7a1rTgZUAe8zJqpGaVRPrZawxs7nImdNOCVmOoPpKVH07aJjjZs
WL7vkusZdQ+jnH7+DDcm8DjllSEcOBKCW3yDdrS6gg4TLBCxZP6Uxw3wtYNWekR5Y1Tk3VXVVY54
9HrsmFi8MMj9Gq1KEjXDqRy1g7ue6jRuZx8Hwv46AflBkRczSX7NkToamusdfqiIB/yIJt+9vEj2
DOxob/iAhzl9xwOfi4nNEYrlv8CdnS0ZxCB6qYLXCaS4B0ujnQQB3n1RJR9Bj4l3jMpNlPluetwt
TLokYC5q7lVhhYIf3Ilws5nmJ5d6jVDtpCGrynmZP9Q99lJCuwQSdG7JUaAka8oOADnrQDPoTU4V
7/ay6zRq5hZPy0F36KK+ufO+YRU9F04OnFyc0y23c1Xr9VfL3aI5pYVROgu8lAp+lWZ0CF9hmENm
7cjp4akqI8jb9iK7hRvGyheyyG2bMMReABqklpO9Jx/vNGy6qK79gfKwOvBVGRnuHS8JO8ijRmsi
iFofzI52dEYB4aaMJOztjrJ7PwPu06E4qIPyum33WhwolKEigxHjFftzm/qA2SjABT69d9l+QBpr
dSS5DRYm5r89Htf6FzgCfC21rFiFplTvoI3obN6UfOxh8JQGXJn4NSQmq5nqtsOr/sikETbpIjhQ
cPqaY1xdLGEQuejmiZbDc1D4qfbn+wLZAkP1i+9QzMdBY1qO7jHEE8a71WkKT0/Eng+YikWXaWqn
2+ibJebHjEL6/bUVWcZg/OKMtUVf/i69bkD8pJQwiQrFuqfc1O7MP/YuyjFJbJkBHvw4tMV8TkD+
sAx9ZFI64nbJyxmy9JB8U16klpy7eB4l+iAlE1zfXw80HPqhWqMXMiXAjl3LNlKJwONnvi43a4nA
Xnyo63fEQk79+K2q567Xj+X6QjQwOX45QviodI608jhqojVjxf3Ut0rXcRWutVNo9VD6zK4JwaOl
pF+QqX1qSZm5Xjw87amcA30hhOsQ9i3ha0YlAE0hE1qtJzWZzvv/9ty7B4qaIinkfBXShOtPrEp4
ika08/K2H3QOHYHZ/3X5hGFhemHvDOKJjYFoyCMOY5dU24OcNABXGw+5AHHbRKjmRtT8Iazg3uW1
joEWBFG2Xro3vVfUQ1lFPs4qX4eHLEWjyrzG7i1Aq2PDQIZn+ftk3Ugjx9IRDCQ8u3QNQa57uiu9
p8tB+ykvuPZEg33lv5GZq9+39YHk4nsYQiEYRXgwvMQmT7O13J31fqpRYp3Xk5LVFNnuS08jhcvN
q17yWUzpefMBaDqzIJd/lxUcrPr5VAIqj6xXtsmXu3K2rgt0SDZUcAUVcvBEyFaD7ZLifnZRRYOq
4PaMnezpldiBU6jV0f09fV+Wnx09IIXEs0BecKKKF5H4A8cwexP4xZT2XAJnG4sAYth6rhW4TOiB
JL4/Fq3u0Y9Sf/8g0dTRQv5T7FchFeCuFC4uWUcO4jFFZzheWrug3nhjmtkKSSN4WC4PHgbtOxYs
KTlRb5WeYYMI5u1IO0M55ssFApX8EVPkSWuwZxerC3fGTbiHsZaYAtzwQc6cvT4lyyjJHqXpHk89
4DqvMZtFfdrtthZGXBeLXcYkQnUxUD+109bVPImBw/75zEzf0Zx9QMjRLH+DqTl7wv3BbBFFXOch
Ci/CkBzYKsx/doNGXqRWIfkDAo69BE9xh+f/DwNae+t+M/DqY4gqvSN/Tv75WzMIR4IXuZQpITlM
L5NWMbO3YrklC4HhK7vFD44uxFgMTq8bYEnsvFCG04FLQs1bLofTxM95w5hqzAHp8zLvwXi1rl3y
ID2fbD/Ao7xlRvaOogdEUT/JvOjv2biI2VZWoX/IAah2Ou9ehd36VtxqO7FAqdXh2X2mVExE0V4o
mXCh6BqvHCuLRa3P17FQXtEA64h1KXUmvIQUcSgQhrR+F5l0KJ8vdkdj4nPDZQKJPFGLtACU6U5N
OnYFs1VG9CLr8Y1O8ihGc57rpbh+7OSBnYDfFYgzN5+rHxsTMDLHHtIo1Ey6vK9kfBAzE3OrOAMl
8CcrYtA5CAW6gddPoOCTTjv8U4Swe0Kq5QrPGsK8IXybHRoZ7MoMMW8uG1UgctcSFcs8OAuo30b7
+E+UfFkwmY6/pUKdgic9HpgbjpDjL2WX8UcYJgDhws9IAatBsTuiYyJ739RZcz3bQD49WkIdM4uh
OSePTwmgf8EeuF+EJD8xi5p+d9EPDnfVDnXRbRp8b23CJHa8Tl4Q7pMKDTBXYhHtX6mGHnHC9l2x
p2YrT5ghX12aWY/0CPd9H/76sghxrVMgnqkbVBrYI8zBhWv8ju3wJ/EKqeFL8ligswgspLPC8wAg
yHO/yynDN5yORlf+vPnJLmkIDvfjU0gLxeyBhatEPiC88aoGA+w+X/rhqfkv5Zs+zxIqSCNKv8Ju
2n8R0DQWkAcS4Lg6B51RbwGEe+5tAQwYXFo32kE26hztyCtSk8xhdYnYqt/v2bc3Bx/BilZD52JF
TjCaO0E4BOt1LZwa5iwwq7U60P1nWlbmA1hlSieINGC8FVUxR3pf1WimeGY+zpzQbjK2yIehzFnJ
gkVBAhFUDmSG+rUSAUd0gBg34gSgsXsqy9n8PLZHEYIZBHt+umfmNOuKE/JgaPlHJ68tHFKblfyy
FTtctW9E3yJiXMPvgQs5izfk8Ygd0+SsVKmBi09MN4GcCSH2OCeMTShiDSk0djUbO4AVBShG+azr
wLgKU2Tt6F7cTJ4C5IIhBFRohYR0GQg8aoDBd8Ifp9p2Pa/SMuRqxQ0AT4iUseyjfov2bkOR57gy
kdh5YPWW4V/xzaLKd3YYDoF0AJknI5Dqwb4A2HMmb04Zzp5JFh67IrDYVB1DD1JWN1ye4LXrTVFa
6MiWxVQtf8Yk7yLA7wzO/eRnhKLQm9F2VUuL4wZDv1WBub4hraC/XXzLCFQxM3qUL46RFK4mRNjL
EhAMEm/ikCQhBrcrx/C7eqtVHogQ+SaeA82skJYkSNV2O8HpbeKLpBFpGvWohjNmoJ5Y+9E9Fa2k
QkCs+VhnhxIBVXvdy4OQ4zwQVLIH3IfYqk2eXE6U2D4CNQoZZpuW4YFdGSyTJE7ZKSf7QQFU0+sd
QMRKo6WT9KZJs2SF/w3iuNBy6BfgL3nTFKfeeDaDaUW6yfyfbA5hMw7i/tuEBtvCitYi78mw2FcI
owAm5Zjxorw1q52dG0yjcZure/2FKv5ka1UK5shnKIrgZ/LXYUZstZi8qzwIsRdxT7itxo/VxJ3d
8eD86IQnTzuB3oCePUGqFigmNgzGPVmkIworq6GlzUZb8KQV1Ij3WbKQXFA3dLMe6OKt/p88qk40
rzqHiwDKnCDkpXUPdSzBf1QzzQRMJITLu+2x+wrTF+FnQ4UVO4JVMa7yxbQOyiMw5na8xY2Stt8U
sqrjF/jxROx1si+eKSfBPuDH/+pXQQPW3pYkl4tOf1nS1Rmb7s5JP+bjcGwuqKg2p/fxeGwOZC1W
J4owX0Q9D3KIAaaycCwTxI2YOgCbkAxpN+FhuuUxqtUg/MEOlSw3YgRLV9gwdi3Mt3vTws5gLSaD
cb4bL0Z7RP7edN4n40f8+atJTl+0pgEmr4X7Rm4mFZ2k4RPtyIxtVMQr27xVurN66I/dshm9dFC3
8xfIkqd2io4mQwMSQlg6wgJMQTS/TPzGInNcgHjdNtbSElpjhtweQRtZP51D3GTJstu8mwkg1rZG
lJQ69Vn+S6uffc57YPgdsaoP/rTpcGADCl2OC1g/CEiE79VuMCZS7RdVYKYJq0EjTMQfyZ/KzOoV
ygFQvKktjDvLuo6WyiHvQw37MdiaB3ElCT/9ARuLBmMle15WuNxFGmXVeTpo2Qr+q7fHYbG4HlUB
7gRNgfXw1HYqjwiEUcsmOzpU3dw4zOKIipU9qT2zh0Roimk+ReQjxBWIOGevLZn6O4IffjVwrvnA
NlZacZmjwm3saxVMxAOBLv9KvEdAObM1VQizPi3BORcN3udo9RICoV4wywSRWuDO6Ic2RWZUS+2E
cJ8AvNx3ipImZr/QDNaCBX8OdtR6FXh4LHlPJDODMjQEUiiKkNFTB8IcM/TepUQmQC9ouZ2dgdsN
1Pv1Qx42io2wPbH9oRbYWKDlK8+8m/e36G69P9l0fkLP2RRfBg3icNiq9ovS9waCB4QgfC5fQRco
PPQhkVO4KCZeqwKnHQss66FqwRV7ELw+4eIehgW4AYSHWzyArQhOLiLeFUzFaDMlWqIke2avF7jT
d9o8kcDtChYu5i4m6lixXenWP5JQ2JQxNSFZ8V81kNYzQBYdRbqMALm0ITAWkYN0zsQsAEraXCs6
KQJKkRpKwocPfWhyu/NuMlyq/d/+6wSIJV8G4K4lRj2CYx1HOWEHF7J4C+2yD3J+xKfNurbdbih8
rQPnkC91CTH3bO70sDp2doAV/P1MtkodYcmli4cCFJic/+rjf+GMxN8gvYM2w12ZbDEeleF/obfD
oWuNuIpKJWNJbUnqAH/WefK6Kx6JD0u+NPRQnRfQFclYWG9ZL06y4Pz5VZtqC4zyJFKipjw+RNI4
Q/zrCxetqUMpSDVdDpCB76bvYs6kjL3xsb2lfpesyEW25+DadIEP29KKR5BOKxqju68DxW9wDVm1
LasFj/3s5rOB1GRMHcp0DEhM6WlE6holS1EVECnM/3mdntgBvGCncTriLHKCZ/DkgT6fCerUQl4d
2vyYkSa6EFdo3xofjfAhd84ILxM9fZlXtzOTVMyh+GFm/u1r4PdtcAIXfCPXpymW1zU5nV3GNYpo
3eEk2OfxrDWMDMXH3DT9inkYMJpJMonuOlsl0CTxRoXY3SDHzt1Tt2hkCj5ACr5NPalPJ4SnhyX5
GdVSgppG1e9pSSPowFbKfotgF80wyG32kDMQ+2xtad05dI/DXDsi6XuDEhPvK0PGqJrv+1ujlwQg
iNkeVAkfnLm8lKlJR1UfOlB1Fr9a9lmiw3naFNptMuboeARhyTJPzrWB22xh+k1tyFfXUzmvkm9B
Bn9TwHyM70JnYCLk5ybypAHiYp8zhtqdoqMplC3irofAdC01BLEKv7bHR02PhtBQIFqWulxIgrmy
KnkhETsu2WtcwsDdbB1INgE6xurAg3nPVfwFxbiR97fP/USlnwgqRntoxAruuPjbQ9OL8jUgRUVF
vRIpFbH1/M5CmEroT/0UykQyGgwVYl0N6nC16F7maKH4Ejm9zjbieonfQ6GA5lh8hTbIwh1LH5+j
qmqNS/i7WmownDI3sSN+UyX4U219wDxcLDp3Yj/NmWrv/WYsGkJ/ArPDqMkhqzJGu5KEcycek4K1
GDCOu+VhLOEEUXQJrsA8dZRNDN41ZS1sKz059ZqMvjIpSf0emXBM0cZXeplucjqeXzTEJdayF+7M
x7aMTKf4skhy68mp5nli8VOn8zjEIAuy+ISIkgpVj755PDr0wgGH4QQfaXX15Dcz5eRaIj90eMiG
n0NjAIa0nDOZQBj3VgFN3+sZCxmXiIPOZ7pKfPH5tJXlRnkKY4xapdDr0VmfvCdAiVDWm75nnXCF
Tx359/VG9PRiDbRW/frvqKNNxTMo+6lLW07lb0DFmpqrcXnSF95ile7jpOtHv9DdeMFv10bJbPhd
LEzJ+giKFROlXiM2vMr64Qjl1DiQx1DiO8JFGdUY1PLeEiK2rXRe7Tw9jGLJEDZFwhk716a9SGQ7
DQpHRnsLF0Izobf8vFWX8q6iVp1mdUmBKDRTU+2Sgwka85X7nCvl1fGmWLVkIg5SX1DgFxZqdlPp
IaZWqGi/2rxn9h+wuLOQgbLXE9NdHHXT53EdQQcnFNn/S7clL8I6B/cNr9wEgVPa7XvPdX0xPNaq
OQttFLChkX/7QzlMisfzXDGxhOVMX4I9pPDh2kjB+Z46Ym1FeW6eBDjGYjKUd6DdxGY9P8AUfqpR
gxXdRju095dhYFLbTZDt9kI5bJGiDJ56Q5TH6MUjz+tE8iZVMLiyn0fMO2+Uj3SOo+jXsvPI/AJ/
Nty3D4O5P2eT/8JadXQ1iq0czCk2QBvE5pLrEbyHmvksO3UOAoPNjJbZL2BmUhpk8r1qNFqA5PBc
CdbB7vJ29+h2kccdk2FVMzjVWNR3bbasDOUg3YnhFPI1Xw0ZvauqjOAcUq/WTEM3a/2fRkWuiBkc
Qdp/rTrOpFVVA71oOdv8AcJc9lPGdbSm39UBE04jJ1badv3G09vST81yAcgu1pb6ujZ+qVynqSOE
0JJ78Fr8SOJmL07mCNvwQI8FqybIEbOibKoM22bfwpHA23br089oeVzKw0dg13GxLrthcdrra7zs
ZVuXv1pmpWxlRZ3+rHPWCrXdGl7cWjuVJGbybzyx5ckyzlp/HJM6PmFUh6KiDOICLG5TN0WMd/gx
Yj4TWVbElX37Swx35TiwHRIga3rAixrQMBM8YWL8NpSVZvnSHJbadp6j9X4q6ITtd1sAPNwKWIoq
mryAR3ZiwjJpFx6IBiE6ZPb1ZgG8gChXGgA+8jPAH4v4tlQO0/tlq5b9YlAlKlsVAcP9K5jhApI/
Kn0lz/0nwPzWd4glfw/bxXij/9NRnDV4oS12N9vdo2XlPRtxQJ6vHKSgWidu3OhlhgW9iMwS4ocH
PAUOi/goOYeLU2Qn9hNtnUclU3uXzNn5XIlwABxeCTbtNl7RrEzpJwnlTcg/1DOvK9+B0yuDp8mR
6jWWTduxAL2jmG3hrixjy5QtJ4s4CSRKbIdu9uYuSxJN5c+Mf46yn0jrfotTgAp+c6eWQsUSoR9e
Mrh360GKXeLsNsboav15bB3d31TwS/ikotQd1KtiwcWP+JZWBaGObbf9Ym8jhY8nG73YJCX1xEGn
TZsMIHUCm+KIJUUECpyVHRW0YJD06xYQ+7bZVrBYbh9uzBm61YtYzdEK7Xr1rgZyut/V/Pn1zGV/
9a8fwEwl+sUJ8GqZvDKQAyccfyebXWTwGnLpNbz1VuuJi8NH/evnd9j489yR8R9a6cmzIt173b8G
kvLN9pOLQJf7K3TDb/MlVBh2OKDRFMXn6c34KyzTYiLo+gG6aST+5r4Q5aA7c1mN6lppP3mMOdUJ
5cNu4OLIhlwWJJB0+OgyhRwrXX7Ow3Alj3X02an+D3kDp3/gqecxWceDAaO6SORJs8Br3nmi0BXi
G66sAsBkbmvk2vSz/dHX9HKfqoy/r23KMf64d9jDaVJV3clGhJyqZ9TapsP4hKLmNhXfHzWY5pjS
X0itjNRTf3dLOCFgrJg6EMIpXUz4vxCbeIIMH7FQKYtl8U98DN+LT3eFDrSuAYnpkSP8SwoDWs6K
z6zZ+eQk9j65lFnEFOL4CuvQfM5S6lvZ4upzMJ4uWLZLz8RTquAnczpkXoxuQDFHeVrGHHj2Cjax
nt270a4ZaP9db8q3HvRrMK4NKYZ3gViOBudIIHXCLObVEfCxhUKmE6G69h38Kv0TdwEV8fweYiwk
fTjYfaONW1YFDrUFXTLAxyxId98BmAnGZ4SLovWg/oNHu90Nq5YPgjHef7Qr5EclpMBwjJBzFiba
kLu4qhC2EwJpx50cGH5IDbVndSVULB9MBj3MyC0m+s/aRED+BTCaf2q8gGPwzsMmVDgqSTSalMtm
v/o/xE6CGduUolPJum+XYJRy/p6mNrY/4FfYQhoS/5amaW0cIk5A3tIvBAGRqhWb1PD+m/CHw1mq
S+FQcJJIp6Sbt4ChHdsAZ7Awq2jSa95Qemsy77Pw0N0JOlsot5kqiCik6X3dl9yvshfMKu5Hgqhi
WyHSrDzmJ1t+10gSe3pRaQc8WjNVRG1/yozV9HrEZ7OJPCmaqKNRKGMUKDMtNhRnB/+lsXhNRSb1
nJPMNjMIyvZT14MFXnHyahxr/rq2gz541n5Gfq4LuTY8udvsX3pYkm780BuiBh3bI7vfkNzzvNqG
BExz3WNXZuJkHFpm264yX1aEG3zPLJuTxZRzELfZDdhrkh3n6IBmYoh3wv0ZqkGcU32dkrGWbdBq
RNW4m9k1bdMO44/0zaoQTF4dokoVHTyZcQDH3AcNDDvxwtMmCHNja1alOU5Z04LjL6DJHD8z7lty
pCwvcz7JmPqroQPS0faExrvSuq3YDkP7HeopmTV+7uMfkcSScxJUt00IHr/j6rxdvJxlAwjmQ9oS
5UJrFECJmYO8gaHbRZe2OuLjk5znIkH/T8PlQS0TAOEqoCOmWoBCEN57oRNj4G1ca5glG9mUE5bA
H7P0EQHD2+As7z5N6Tf8/lEZSMd4WXosFiKOtUQK3q507/BYfO1bVGQqUoIZWG9Qem82+vbIzZWO
EPy0wrkPJIAmBYKAkDd3YPB0GkAroE+FmWpK2BXTdGVk7XYYGYeKJmz7UFRV8hb9eXBmjZ3tE6sy
07DPZD3NR0yKroIij2zxxE8wlzATrVZ4Sobipe1+05pQdeoHsqjLDEfDEiEtlpL910FYR+AmyLJZ
oTFV1D+llKSK9zXmdbOgURVfVByQ+sYMbqT7THt8BI53a/15icj1tFXbxsO+Q46BtcccEIWaNtgT
yOoZp2Yi1ScJVoGCHrt7XyjhN8HCJQ4DR2fmyHgZhslXTjXTxYMTsXzLGYMdfIa1ASrU99hO2kRk
Hv1MXip9CQzxhAZkmzNEPvuLrZ2ktiqGEA+bGLifYCbij1ICIaHdA0H6bSbc3QKfPg1KjmUNomCX
q8aFJPblsOLcCoKXfwPifFgLgnMnrh4DNHn8Ovin1IokkFwtcjV9z6RkcD4nHqiErh1FsHxI2fk2
QVUUF6/MqaR7Su+LfFrtSEwNOM8YzxuSMLFfEyhJmKNdmjhqg6WDeC4kIAbHLlhv4Eml5r1MfxaC
y+Rn4iNWjFLLRfDlVextXwW4Ff5+8khwU003H6cBBC3Lp2GtO7fnbfIUVRHnEZhjtjcegHhAarIY
hd25Nj3pfx9zwyLpfz+RK+3xW9k6uZh5RKG4oJtIctxqeq/PFsnHxCnJmkfRtUNqDoprtvAYM1GW
M5Ox4J5E2deVNCmqIyfkxpABMS0IM3CqZGmxcwYQ27tHGXwlXCUK6rkME7Eb8I6BZFjndb5GlOeQ
3GtZhckywjdEYCBXaaxQfILB0aM/+5J8c0WPHKsmktGm295I/UkKS3JqTmga8OtxlAjjzkj3QJNj
Kkl5SYsNSo5Fmdq7wLj5DrrWRX3hg3FP/xcEbSTwLSxOcOqnVzUvfVsXHJgfgVFHB167gbcMUYGv
Ij/Ircv1H0BNglS1soJ4IUpIRLnxIzDxN9UKK2+sDOAIUJdysBKPvMRedeGTO5pICbtmTaik4j3D
D/282Qn1fOr2nPyWq1ovmf5exdaKCR2Aqag/qDzaOLvWY/zKSzs4mJkfkaqOC7o2El3Dra3n79W8
I6yfmL0Vjx/4RXmmgQh6oL3S1Qj/uyRjF2+qEJ1Xy2+rFFSkPEbQMOMULK6L8qj32585hT//ArxU
WeXp8OM3VQ64CGuGJ49soLVrk3L0Hx5x4Dt6FAurZdtz4bLEDaWhbYlZonNGHICuyxmAK2a95v9i
pJ+0xvGhiL/+kGIvBXxItqVPF8I7dqFg20BqSOvocPSjB8MnnxEqG5kGV1AaSU/T2eOLvS6IxcKS
/g8K3Hylh8bFpM4oYlxIGQ5OJzmQ9OCDEnd5wSg+O9HosBpwZ1dHex5CW7EmeXb1WBnUi/pqyXxK
x1aIdEfcYxchgSmhgpGw0e17vaxqd8C2AgpDdjf+MvRPGzSUHxg0JnLPdMeE6iy/qHg8oYcftNT4
5uPY0XRLQISXsd2FaRV64otz9taXOUsOHFrsxfH5WCuJ9FDHdM+dP7ykES+ocJse/+KdpB5iKEYQ
3st3Q8DprbwOE3cUOdKAuGk6uru+rQnO9uCZ9LQpK143DN14mqB1DfI+6LRy0D4l6ydknU7B3S1i
lHFSiOrK83bkXvbbOKXOUw3QtBIKIUPvs3nqOZC4x+5ZXhIBqZ3QWLfXXUJls4m3Dbyk/vob1MlM
0In3584+J96CoGnwwcR9dOCcZIO8emP+OsIAYdA4XOQIxssMt30wfsOEoOLqUo6x5L2KKr11Q6uN
asSq9GUqbzM0KHDS+Mmglp/IFyD/GYvGoT99Kqhc9pS0F27rbDyH79dss8M2KYGm9JMyrgqFZ2k0
5vW8Pu1OwwOaXhRcwIvZtmPW774UhkXVU3LF0E+Jd4elmg1d0KVq2YkoffgelLw1/tCooH7bVwmB
NbGSHgKrg2GeWqlG/5lvNfgKoA8T6v0somfWof3GTCsZaGeq+FduJAucaajm4xUq8O/O28M41kh6
iunw1yKJaDe/CrM+TqctmvCX/uhlEqQFGdhnJEDHidVF+UlfVbIY8tbYVbAGy6CbrITFicqvxSXY
rxwVmm4s5IQqk+oo3WV/tON7X2++MMZaXdTF5rZmmqU1Y2t2vzIWzWQqBuanvBgKjQN30j+aztde
Yb5FsaD0MmIZCSfAP1N35GQqAc4HlpTjiog8Bx83NoDpx/PtRWP9SzZmQgfg5qrbSZqs82MmZCjo
0tvKU56/+ZFLXWVXgPqpGp8W3GmY99RLV5r6Z97ZNn5NCq6qFiSprde3SNXjJpuGyohxp9b+x3EP
j+oaOSWxjxp41//Q6hJ2EXJqqX6rM5bp/5w9zc39yNCmZibYcUC9b9CYkB+wSpM+r4x4mbXOGpSv
cqpxxWtTN/iJtEJolOnLGutrHpVTWR+hMH+01lVVqIksOYqiGt7OvsnEdczBD5FsbtSQRJRgw8QS
vSxU4/onoxzP6mL1nIQkpyYrLBOxXC5HV3ou7PVxCKYp92LWw1UqsS/CUN8zB8QJywJdSakEXTz5
reQZmynaMNUeLg6ecKxRkW/VuttDUme5H35VhYjCtCG0/SPUW8OlVunufTvKudJZtLJ4bzWjPo03
iP1S0JwS48CUXFMO3LV1rf9YH1CJxGvVnU1o42tbsCGFnK/J5UyhsxFeQCYeQBPCByzWly1k/vO1
1+HUrrJ3dplsr/fv/9/QCPaVCFdMvH02jWDRt4jdzLMA0AsIXgct4sZLKzEL7EwCoHO+kYnkJmNP
du7xJXWkiRHs+Ut+ZKLWSSUJ1R6SM/jbZ370GKQlLriY6sBHUG8aHzdMIZMxsNewsDgPlKiru6bB
qKpFtur2VL0+w6rSrwPhR58MSfcYPDQiBwOqrRocGkOwk3rmoxf0H7P9YDe6m/IRNVi4FhcoVc1h
l3IVAi+10+F5apbGiT2jkfBDz/u8DeNND3RSbLoihtd0uAvVKjJENVtr60REx99YkVcEcKWbBYM/
Fvw8p+oR/1Peqamz6cLuciZBOjI/FXNz+nugVdvr/zO+vA4KLZH7oFzX6QqAT9u407X41c0uCt89
N9wDOoQbFBdRWerIYU1XVOXD2DUhtkdA4U8aTy4l0RGOaIf8goa8oam9fFi2IyPav+6j5Cu60kvL
+dgV+ulIksEmZ+Ya2zxfTxD5oo/ZVBhRzEaRulDSlGQK6g5/D8qCjIsgaz/OQqNvt1a8llJHDF6o
Wii+I5mExH4EVLVb7ItA3+RBiH+rK4R4132pnHMdwbVQ2FTqttV3rTRP9u25z7T5D26M8lzOar16
1EakE6om6CFkI/Lk2duHH5cXFSdg2iHbGuwjwkKRDcPjoYYbwOst1dL+LKLZBeWmzUBdg9ShQFr7
4OZUs8dBG3z5qhROQyPaa9kSI19q7ppHPyornG/6lwemaPDH8kSzS5DcUgItbMPTQdo5pMa00Pr5
c2G/0yOADz9n3qCdxiYxMoSG5yRM02JSWxJGVsClOWbw/vjs5NNGvaICMN4CbICpfcAtdzpPPAdf
YziOl+Z7V8XotbkBCdVsP9xoOUpQ25uejcx6AzjbvVcZrVuODym339qYzGkV99mrNujud416voyx
E293UTDHsaSIFbvmGU/oLJzpP0eiDKMtr1lDElYh/K+S4tjc3fA1PZX2UDctGutcGY0BjnfQheMq
1cA0lZbhp6Ihw5rPhnF6Uwu6af6dZQAetPY6yxlVZPaqaVF1Wx7O6CCPKgXwxQCC9KuoRpAA6+e7
UPBDYtzFNVT+/8m1bOZwLipbnFMYv/IdKSpV9QJrMOHI9/wIUldrwuISE8HtGkYYe80HTs8VQOq4
zfipIk4kXM69ofKT3DckeK58YyAR9X5Rilydm/W+7m+Iz55NxKSd992PjAEEeT1/eRa9JeZk/iWu
THGz7OusImjbR72jDTYH38V+eq0NnOxlzILmi80hdK0nm848EUBb6Lvg4fNy+hdH2VdkvyUmGO1X
csIA9FZTn6w1FeJwQARyf2q912NLpa243oRVmL7iKroViM+3VcG9UrPW5zhtktoCOF85E4Z6XJm8
2wdD6fKXCVUiclAQfoFOJgp5jfGyIrLnv/ZR6psvmBFpK8WVoQnjqv3eyTFGBaGU+CEUl3z+y4lH
glsfw/EtmCY5pwjewNVyo+RjbtrTQV2D5FRvY84HLlRcIrvTnFgLnQoCbDbpwtslhVKgGVD8CdjU
ib626qtXbipveGe30fKuOEEn7pLByEbmGOQHGuO/rzpuiBaGFUppAKvIespkhjnpa6065DQPlvvg
zJ9wpzYa4/QeqzxIth3m5cc9kfhGopJBj1X/TpUPpx91bLZQUK5hcXJO8V1XTf5sa+67KixmRgrG
A1uBLwE4CDywFMk9apdKK7x6h6We4eqrBRmUU3FmQXYe0IY6GHjZ78ktjP9SHOYjfRV3/Hto2z69
Qbkw2VsnumRvRggIZiqpxPpqO3HjmKbXBgqGnrc4Gjv+2tPSR/gL+i2ClfSzJhBQhMIoM918rV5c
Pz9dTca9LAqxCtxpnMjDmidgIIEL2KrQeitAYWwliQ56Ctb2Zx0KE3UJW53A2YGIjovL7eT7//4R
gFEbMZTisW/EfcUTdL9wbvEfUcN9JhatZZ5Gm5MzlUl28MLGB6s5AfyDUNS0WuwBS8lSgRUuxNpP
NnGyMWtxpXQMxPgW1tUnjdNuiAtCD9amVfTqPYLfYwrayg7f59Ku0/DmSR7GEOzXREtcAox+HA7A
3eftW0pQjKFX0lnjwI8iNj149cVdm1AuQ178Dcv/gtM8ZAMQOdIEqbl6kpxZVXUrf2MkbjnOSRu7
mrQI0IVfeXE0e+AALiynrWmMEFqnJQzfWjj17evI0VCwlgn8g0DF9QrfuR14/FNVjkxh/rpCTVb+
cHzxsJKJbSQauznPEZDAnjSAPv2ejbnYJhc0v9f7WHIpTbiNzYQlkNlJt/PpzOpjI2kpQ6He+WQQ
MAyJkicOSyiafOwD1MRJg9Ivdv4g8ZXPbLlFH6Ey7gSwFCm99K0zvpmZwSWRVjMLSBWscxaarkrm
gPN4rfXpUit0thr5lnzRLT8lYFUjHC0WTYPmr6XABiG8e++qULpg2mXQ+uDnB1+UMqebKqkcu4tI
BvQpyCFsKFT2zKEvQS362tcjI9zS9YZ3k9upyEBgMkrFqAssBweewsLmIjIfN99LvMvVjC8kc9Yz
3o4WboopnTdud5DMw+wRKR0+x7zNC9VD4lW1Yqh22cYIGxutW4/gAjJgXeIWBdIvO1hvhOekH0GC
lrcKWEiEt3BJkmq2c83DCCTn0JkvUy69vq7CX0oqYsqWfT43zmdhW+7yIP90I2JeyefNYVusWWpg
0PGPau7fL/Rrd9q0ar5Eifq3SeySTdOqtvW4NPeMS7pTzNw7Isdg9sz9y8vrXbct87AGSBeVpm1d
kxdtfeQeL5CTMaudmM9ZoGSXPIel8mVY3YqDyDa557VBTd4kErNfThanMvVEyWNRjVhirDup2yCM
rvvZu2AD0wFv6gT7ym6/PAj8jNAtfltEkaVa/AuTWplbcmocwAurONkSOE3bZR8sG59M/+shQEHz
h7AL7fUw0tuuhoyOfqlwZWsaFhUO1BICZsUUrexvKiNKwCV4y7y038Bzxc/y+c8Rd57xkzgoVID5
PRzXgCgODxVB5TdKa6iVC8h0CZmPsVcoI1x8ZgLL+0KlFqcOEKdcGYhuwRwr7DhpihneYW5QDgDT
4KmhrpmI+ngE6nPlZxd3m11YEufo1ZZjETW53/KRKzkVFVnfzympYZGw6atBOCPtQKC5Wy8GIFn9
ZTTfgIUu95AUw8KX0TNsbxF9QjWmuMg4O3EeeuQ7fYmKqs36PD0iJxNi8qNH17tdKLuxEbIppZwh
CZoD5ZyPbyk+8wxp6xlpmz9JVJYsf8V0lc7WS0ZU/GSJv90tYtapWEAGdl2IjK0VgysHWm6NfhiX
RKzhWzUb8Ll6w2VkDmSAfyqB0bAbZ2PVb4J8TF0eE/PmEuWdd44Y4VRz7KKvI5v2gdIOKjTtZDXy
Fmd5F8dxdcfaAIx+hG1sEsmlIMB+gk3aVlrslc6AAVbr+7viiHecupN6XvIMSyEAv3z0Hhv1FtCl
T6FSRKtL1ulcQI0koj+oYo4L2WWpq6HRYYvVvrluPVLrBXy9V4VgsF0ZoTh7Fm7lbXomXDd9lCL1
exbAuhYT4y3em6JjUH8d00j6uY1frg6o0dPRz2fRMgN7e7oixyFeQFNgN+O1Etv9HSNrpojpwi3o
MccXFcHnbqn7Y7J3FKTcZC7rPCvfwEghzglzud38KOJaNXnZ6fx9L6lcxhi+FNSaxHY6vyN6y0IE
wSBAss0ZXTFBvlO7sFkIGZyuNTGDmzzCwGsnV1zpRs48fWcC/cV1V+opeVey1+qyx6euefHLo25l
7R2dU+eLZjIZfuOrDGx5NjEILNlRsQ5VUDPy+cCkH5Zc9H+8o7K64BncYX3qjTQVT1bciNcXRaAs
cxi74w4m1EG/hnCF92PCsXbzKMDb6UCODU84wtjJ3S6pHV2UNWChaAxoPl93aF9NhpTj5SsDL2Z0
BMjO2IhkesmSVWKNPIKtIqthj+cFUXWbgqWSpoGCe1vyOhuYQzBm8S0vhfc/PdJ+4ujb3JuMXEVU
iy6T/OwjnyeHSz6jmev5Qd9cqyE926+r7Yl2XgYklgti+CX6PKYXXJI4HS571Wb6eOZ8Y1b3C+Y9
0ukfvCzbd8k3qT3LW6lz+nHKspHhM/C0PX/5vudRn/2MB9IoRuyLIaHvKlOWRZ/4oxBps3GrVnnS
wU0+31VJapdeCaJBGpOJ+qqg7w3E6FuM0h9h2fJsyMjCr90x42JDkzlEwm77uepuWHZ1DjHpmsLc
Get5NSs2lYIaqkXx14+2bDE6n0oIeqbSvHSbbvE8EROrCQsgxMkx0I4I3OO0xWopct1hc01J/eka
Mb0ePmAkLX90imdB6h3j5stu2TCIPyIVsObAGsOvB76p6DlcTsS/Rr3LEPKQtVJopuFFJ1x+XszL
GiUAMg8uV2B+tevqu/EcgJFNHuiKRD08Toul4MxhqGnbIPwSl7p1wW6xbLR9RYN/7YUe5JXXvrf5
YA95hwTKjvDS9KYqAiU821balbzIubyi/FIgwmVhJ6uYRRiezQHpFbkEMA5HmS13Eb7CH2Jclhdp
HwBTDbZAN4rhCX1bWtQOHSUoU+PuA+TqMR46IBwD8dwRs/C6PjijoyV6IlPQhN0sOAQuza0bNlIE
Z81M4GHWIY70fRXE3L+FgGIE1KJbRuB6uEC4jXYW/gk0e2IHxjVbCFZUfYVMZyQn9FpextIe+5Fn
wQmNmEPFzkkHLi1ACe+N/fqtWLxt2JOmXP0UKNUSWhIkamybVHL31fpe2+3EjarvWPGlnVWG39y9
JvbHL5B08oXBMp06wdUfYqXbukobbRlw0l2U6L7UWBTxPUNzO4FmOqtkM1sR/kH8YSGCIM/v2bot
rS1URSRPixEbURpixoCwunW8mS8UQ9uSHQ7+sZ2aMA2zDIKEJpN2/V5rw4JqdJ3CU4B2zW5Qx9De
LFSVeMeqFMNtv3Z+3ihkvTR7N9CFO5ZDBirYEAkz5k6fMZwgTz/x0H/+/Iwt//4C5PF4A/gjXdmb
es+nHz1HwFFkZtGqVSsFtMw/YPfTPOyZAnb7hvmEwbK2ubMeDdKjTmR3KCKn8oPgclvBWXYytOpE
lXahYFOg8oCnBVoItfIIl+c+VIFUQRWTyexozjp/Z9xLYkkWSjpqjH/TLJIHi050X+bUt3KRT/AI
NFmywD9dGdF6jJlkQCCkZ8BkepcR49gqcOOq8WTJI/DDiIZtOsmDKtfpmybL/026jOHMH2KhuyFJ
f+OhKIPk/DLoJFLG84szW9FxRBHwXJRXKtxX+I43tBJN8PYc19r6fN2pTdQgpqwOIarKYerQGwNY
Gs6w7EYrSHd1mfRQwN5rl0nHm/TrXOPSKXAjzlkL1xfsID6roBKSlbUs0MP7XnwqMXvD+9D/nvZq
xL5DW8auqPDD5OzJRUtrqHcbk3dqOrG+VXkVJnCYJjs21I0kBp0tCVPsWzXghdzQ60Qx+/7+1Oxi
Cktc6jLEf/VektE4cpm/TTYrL/D+wslS3UQm/O8ivG+wDIN4oSWl+NJ8VYi/yo1gin5XzzI5ccDe
/Yid9VZZRAlVF4Zo9DnyaPabRUWJ7l6qO0f/0lKUcllM50DlP75BtkJELZ8bLiz9D1ezxGauMetj
lSdRdaYFyuqeWorebbFyn2/VPFUaw6/WG2uLcs0sIoMsFBkpFXffz8LjjJjaW/WkCSd2dwrEGEZd
upCtsxmfpgZ85QmvTz05DdpUNWPIhT30d3aGAyJi4ijutW5je4I5a78xP/HVqq42Q5muOnQhLNAV
h2N3q94APX25pad7mMrXKwEV5Vd4h2SRGdTpb7D+Pnpc1BEwybDguUfic6qiyalFblxcU7IpLze9
erKI2Zkla0CjbQypeyyH/yWNFFUkEFnnkuXdgOdKKOCEXLUbwZvbj5zcpuvZ568qgbzQQT2tTjNu
K0PKq9yCvJTAR4YXt5tW/Zem8XyUnNAoce5BdffT/Nu74NwthKsi7UEJEO0A+k202sCsJ4QGa534
W1EMsXH2kWXOGv7wbElV39Qq3qWRdgtVSssHrg9oZUDVggvxvfcZslQ2sd7kHakpbTmhqiDE8G+O
BEbBkN5s+b+o5MugYz7bszbxdJ6RbUNZgQcn+dEiik/bojj9+v+p8Nlf7MbrLDNvtmNXFIAD/VHe
fF4efQ1Qfr+XLJZzqO/YS/V+XWWaWExwkp6CiG55967rx0ywUv4EPkKCmX+KAO3a+nUQm5zx6UtW
+4Qw0UljM+6gZO5qvlo+D5HdIK/dU8PoBndlLIoj3Em0Dsfh/Nx257LjMxfKHorreoUIZecq4sue
SmpGCxdB4/ElBDQPXbjtzg3FFrUtr8vEeMPWz3RMbQEHrKhv2g6ZjDmqEObObP+d8wQI4bZq1Y6g
pSye7WBEoO04K4XJ5jLWDWS9tYd9ciNSQQb2ip9V1w7jlEalsSJhbsIWuiJA9XWM5bMwPIXPr0s/
jJTqOppbLj0cXuLWGCLP7O2SAmW9Sg9D0+7BYa5/ryAIVlBAMVKq/uS+FZvbspKJXwQaAsZXexGY
hCfx49nLBEzCHi6vmByNSlnx+pPXGzu9IARN/Cxyn71YYf5BlLNC6/icn8hubO1UVGO60V0kZb8B
24zRxyMxiIYFsLfxnDGQ+CosnQfRK/y1n5omKGhVOvrBfXqewZLZ1N/o5hjXeQx8EkCjO51C9wem
PTRgpijvQioP2tdc4M5N2rI/Cw9Fcz+AnKN5lbt4D31XCQh7SqO6gtySadJzJtq7HKpBSjF+HSZG
2JVBSK9U4+dSIa1TO2sVVhu2FEqG8j88wW/FQSa0cpdbt8LpOoC1tkH1CzqK0KwHjfQ0WpwCp8B9
NTjA2nOipVJ6UDG3sg6B3ILCdyKDEkp0DVH4o0sAUKnSE4CkWQdzeD6+3HFKjS9dxyKwVObTKk2C
5kZHDFkErZ5nS7pFuqVnZqtFmP3jR24FySvNWO3KELllyU1hm+MOkg31mbg15s9lygHajIwTN5a9
3GnYDaEgpG1mu1e9LY5W6FU/nn7Ovx8MLSfdMKpKYJDRY+y70W58k2y/n7xxb+Hfy3rqMaCgGOwz
fZi7pIFZCqocp6oNasVaK3NuFnq0N0kdbHXKrc8OBd8ec1I2mmbpSJui1CeEHE1IVh/83Sex5st+
uqcGzCBDYy6C2ftU3rJJMsJANsues5NFLCKxuvfneDzPOTo+tRqWaZYpZAy7GFVysxpfSQqwr1eT
PKNHPliZ/pqZZ7CRkOkl6c4B2h2hG7wsVeLOFTMkPkRgZ1rnkydAQI76vr54MyRj2O5tzlEIW0Rv
KBFnu0LGGvyBMDD/Xg7xxylo4TcmSYCUqdQtberYTwFPyjw6JNNKOBa3lGX7LvLtQd0seNruVwYR
e/nS/iGzEwi43+3wFBZ0xkz8w3nS1gGqjHpFauS9jA7JlM7nxWm5hJjIZOZOyv/334jtiWSXV6YH
ryOYcXthGH3BJZ/mg6gy8Gh1NO7uOQko8q6lAGuoXClpzcWC2wh0PoXbIo65HAMltIK/VYxlR3dx
qxm8quShA/Nu2+6ZdVY8Zv55s6wbIrENA2rSUvl1ixVANxhr4/fc/CZKU9fDrmcHapfObnRg64VI
G4rvifJAJ08NWDVT8J8OPMTJEamFjSb9j5RO+s6nDMgEd39Tgrnbj5gyKK6cdEBMvnDNqlPbHyzV
4KErvOuzuXT6JEXaB+39tI2cGXZhBBjmE8z4JVR966iVR47Ejj0aqJGxvVmSmZzsY8cdziOv0ZnH
VUR1v0nG3n24OmslXvdev1VV7A7LL+DqCK4ymEj+K4MEdJzOHwUxNIIpHps/vQsqZKFPioW+RkNO
16DOhs7oa3KnNqg71tZjfjAT1SEVqwQK1gaaz17lsEiS/t7kOS358a93635a6Y58MEbQXpyyP6VP
hOiI8iBV7TBg8Na4VvWfBP3zeDzivpZgp9DQ6q6DOZU4jkVOK5vlb0a0jyRb+msQaA1ap4XyD0uv
JUbZfF7nljJxAC3T/Zd6gfzeOm/NOckFL8MzA25x5jvY2ztCJIA/k5/Nh+wBFc2MA24TmV4JrptQ
o9SBzVtXkK82U15Erw7yDluHhFvSl81M+htkvt8fn5HMJ5uof3nJIWomjivjaa8Kjfq+5Ynw7zbQ
mBtPf2AdPaLPO9V6O1+Uj5H9PXED7DkJgQ3dl34NRrHamvm33gShBzMpjCrmrGOpqUFESOYZ0pbb
L3cuN9jYpC6P2L71BIVIiGro28tfSuWuFdXaC+9Jn+9IjNOcnkw0qODsa6wI635hxKv+x2Rnc5Cw
pH4tfKFKWkSct0uBaEhl5+ttFkoTSv+5NF5is2vwgYx/iwD23h0G/9FjrsOCAVu4l2paL/TcJwJm
RteW42HkdnJk8pmJkq3w80Bx4pDzzUcXOFrrhthiYbb8/3RqeZJrN+Rd3SDrEc0XQnBXpAiOIpQW
EE8SWfrdb4olZ2orZ+wcCA8AnN2lAItMSyKRZfmswTUylRF7uV7h3XpB05S7OjI4H9Xfyx6wMMXB
Tb2XTHPgl6yEfuLflfz9xyYUGZlELkmheZx9esyFeoA5yPsEDppUdEdSvePW4PPLvkxpBiq2CY93
Z8uay8BD+OIay3PbQkLW8qf5V2JePAdS61R6rs6EdSBUYjzZKpX5UFgjfFt58vzHFvGVXLrkWuZF
+dCBIvEN7ZKoXtPTo+JDT+CVtu1BhtTqe5BWxWHcsGI3dFCcG43sOvXHvpkQ7Q0KYm6A1m5AN+Ak
lc1WDbfcqR3FLuSVAQsdwD2I8WxpcV0duhmv/QMTZslak07/xrQ28nvdY/e7O++jK6nGrntTUuuQ
nQZMTWH4g2YGhUM51pus8+6AByMvYZPmlAWhDNEks7yNXyMjmklb46JQxeqvY5Gn/Kl/KPk6IAyT
MKd4FFrZY7arzqN5hVfbYP3J8NaEZ0InPH7bWIjAX4xMlyFEPMW/iaN4YWMOv4HKEiijEIv1ydNf
vR5wMHbN6oTLR60uEYiPpEDHECD6zC+paR96idmrLTwU8x35DcfcTMYpkwSrEW5rt8n/5m9fEdjs
pM8ohMQfk/8favwPYCNh+4skvH2FvMEt+KccuBlW92rlPUd96mobbaoTvJ2b5aPILwMKWDiIPYEQ
wAcyljABE7k82k3DAVcLtoMXUj7oQfMqYWhW8ElXX1rFcjeADZ4obUQUz7fJaPOR1bGKIgtr4Zdg
gH8nIf5OL58xuBogDg1mIdFGqrNW7gT1AeVAEl3o1rbpSOQLeTjiGH+KLE2QjwXUKDHpmzX1RDDr
Pjk0P+5Y9wiHyQnQC2CddGwT/GKFJELWop4siWR690bf2lWKVY3/l+jaO7m+w+39+CXCVZncuCqd
RTZkiyCCWFRTwMfB2HCz3rmnTyDvppXOZY54J1ebjAM6Ru6VGzAstuk8ocTTVzoO9LIVKE8/GvIA
ThYt34ACALAB3fafSWvPw2RRlj6lZigHLsO1ew1QuqjwKVtJjD2yeHEkkupDwtyRF62D+sv8S0WJ
OVFC9t72hR3OiHOakaUiuIvR8/qjsqI7lpnSV0XgAyPRSnWN57Pd/emNiL3eHE4CZkr4ovQUqoP1
b8VV2J6kdkS5u1kuJWiAlFlIzTl4/3h/wPSFA7Cm7Z+q2aezh5y3i5pK1sz41/bSObvadpB90IpB
BrTxfjUmptaLpNJGE1lT1qiwHXvh8us14gh9FK3OXmcIRWHxvOOSu4zksZbu/VFCJsEoHmR1qcZ5
+55vDAwsp9/RUe2Dl/b54xhJ7ZKMPVAYmARNle4l2JS1g+SWtb1Onfg/RKHz22YHfTPD2g1MlOb6
Mswq0yZjUwio34pz8Jx6YLI247DZY9nusNmvh32UbzTRG3ux93zaWbrKL+HV+gfCE89D7LFugytT
BIoWIyMZLiUKpto7sOZ47cWlMnIAiya5dLkdC1tGA8p48ZRBcNMVXkfXXz+k7++KO3VyNiQeeUlO
C1AdTjNtCKntxQ30chio8VOZsRuk4Iapby3uTJM8ywf18fsAf+vV+pORfUJ8RYoN5UUlUdxc1Hyx
Jcysl+2i1yDOIB4xsd+iCpl8UQiixC8S6ySvqweQgXHHIb1ZLhTLmoFu0aVpRHMCv0gLnYSztgDs
Uz2mPoaRrKsnXLOEtzVf+cvXfr3KHRZFv7yrgBKTGqv+plJN+HtXXnxFJG38WgexA0RBdiDgGTUU
RuU3sFFuZWjrrqagmcAD6HPdB6uVwLhXZXoyOksH4tf4x39AyMFAO9j43VBVM4W4AvUP/VP4iQdG
9jugFtQKfuTVeSIPmlsDxgwGbg6QAyQ8p0JmAVM0B4iU7rVmCvfEj5vRptOObxpncW5MW7x9ekod
nI4vyXJqXF73mFeOWpKlSBvPtgxX1qK8DF7+MA5o6hqWD/nqfn311+v9G/WxlaPRPtAkq3/MZtcy
edTihjV8/nabcnKPOB2SMvIaVR/msdQioV2jfKB/57Gcz2ck7a38nvHcFus0Vz8/SfKZHRBwup4l
t443ZC9Gm/9+sq/ucTXaR9Ex1PAs76QyoSvshMXnGrOa2FSHGNAJ6uHaiXsgyX6hU8ryKyJcTA9n
HxC/mCC292+iC3iZAsBRNLgLjT0qxfBJSielbsQ2ob/VXSIwd0njjsDOfMSsRLpEwtJ6KEJ6paI+
ebnUbww9CWa8ggBeVsfKaEjTFeyEeYu8+FzsLCKz8rpdp8L7wMtDTnErylfGVJXe1cQ0FdI2S+RQ
Dzx0MWoJp19Uu6QoSpDD7wk+RvU+CVpbwbn3swCMWk7q8NsOT4OtMPBFs5XXOjTiOK0dk7Hpaixa
3eN5uM1lgDnZRtX8U03/5SQw4WnPWrYpA+V2XibtajzCwcOkmKUcgqa1VV4iyQZJ+bs8KyDz8L6U
bTkvV9wczfP8nD4br6UMaOf4l3h6X4lBBqjYbk9z1AfjAiGJ8E0pMJASuz0cDMuRwaMql/32EWKv
XSl4KMNByv4l/pNK2UuRR9uJuL+CWXxAICmIyjvgyg0ob7nEfnuVpd9uxRO5EJ1hzZu+SikNPgqr
BziWPeN1q3fy4Ciq+EmOhKWSAGzcrYIW/eTMG8U+UTp5OMz0pAcHQTtH/+YWeuVEQH6Psx4uvOOw
2pUBssbteFyxc5sIC03JsmKCZWaj8xOluG7oJoJOAbLWmmmk9RQaU+Li4Psp6xG6ja6TkY9+CaVO
HPGi81+CP7o16jaAH+xmQLY3qpxn7RG5e2mX0ndDLKchcMqHtuBaN332vArXYVGSn59AQffQHAwS
gFgTKDGbK5rR5SVQxw0c/Ix6QirNEEvibiTbdcQOYV3X4+M4JC8cpQi7PXZ/ZaeOu4Jop7phR+nk
GYMVTx2X0XuJIIA8o2hARnD8t4T0aTYS82dP8ZbVJX0bRfMVJ8Yx+Hk6xwqwLobWxoJpuRWYDKTd
OaZJSxJxpbWveqJHIqMDCIKMwbf9Q3oESbRhhX1NqZfZZU5fTBbAUaUtZjygKBiSBbfKs9n6pqGS
lfgfYZdsmnKqoS/79NMmqApIZgsMMFk7jFNT+rSGEBxkAclq971UhrbhpCPlHc+XRd+Ynq+KmNig
WBi3qykshRUjCCD0wKqH5QMab7OnDolxcVBCQKSTksC1gVSDZt8YzQLPcsXwMgAORa22vEez7wWv
lb2tvMSphNh1ZrLP1MUjj7nXBDhfvQkPtigtU1n5yv37Qhn96LasZi/5VwnC3mILGqTft4x8kFTA
nxwXHxd8HUJ4AoxXDHwxVAVD+JQpuOQSd8Ei7zhkzOZs/Dk/ty/zP42ip6AQ0/lmQsNoT0e8gCc1
KRn1rw4+sYBKL9K9GXosSq3i6H2JzVv1hB9RQzkkZWNn17rT72XbbA6r1+DM7iSNoh6zg/ZsSgPc
9QrocMOs8LgyivLHbqij3KRtWETijcDyHJXz+FpqNhag201M4aEKoWH+E755IhOeJlbHRSS8O+og
sT1FjxfTNV6vxFMBvrvXSAHsSCGa8akLyPPl4MdTNI6nCsKLwyl8ry7Nd8FY7vX1mHvo8gDFAV2O
QAV1PCI7m7wWqHJj+NK6hVdG+mo0VynBcFQr3SEQZCsRlS2H4bRBw2c3rKa8AefoPoN8UkwlzYtu
VWhjlFMLsLu9TKCVcnLam/7Og2fidiAnHkaCZNECmuIDFTNZxw+OH9yR63xM5ARns/G/A+zl8XpS
L1EiuW7VWY7vuo/qj+sx6bL0ThVUePqmUz5Bir1xvnwbPMv/+3ret227odLoOgBGjRy3DJhYYLfT
pfx9tVHuIERqdUgsp5XshFNG0yiZomBPYU1erTqnThfXHICGQe8pDh/ezL9Z8n1XS7OiA15o9DD0
4Np7hucV9NcanLb7H3G90cN2IhkxkecXf4T8G/8rqSCUFRVnU1FbffFxXaaJHLtvz6kK4qLX/YBp
UVOETeQ5y0JgUhlvrgFDyETGJ5/ETRWZ+mymSAXlcL8hIqr5c69NF4865MIETbnAFB3xAQM91JdH
/J04HwgkxeFQf4M5X7xDHSo8+j4fQHFZTCwpm9tZWp4ClV4cbePbcoJNpUJGklSQFoybfp4ShiLq
P3aEnLvBv1v9tSllb9WnzP12Dew4DR3iN34tJPgxNpAIsT+t0Y39BgmntCWyu9Cx83F72609rJbk
qQNr7I2qW1gRv18qEEPi+s89IvBg74pxeZx73pzUzG/CW42EsFzRa5D3Bbyo8oZRCY2v9qxsQyi5
AuxwJe2O7dJUC96SldeJ2kt6M9w+zMSpAaDNDRn+9HVVDOiHzfvTK1h595Fwo9xKxaQNX/UOWNO1
VBbLYQwrv8jPEA2aGdCZrbkGLYKKTXwFrbnFmGmizqHONfojFj4csU6IEsbQyrOOt5sTvA5qg8xL
/HFH/UmNoQq3KMa46D9nlBiu1aSCkfhxXODRAwpbmWzhkBRYrgI1fsB2pyf92ebqROuCXMMCIISd
GdWrhoJKfGSriznKZM12cKuwyPi3SA3T4NjkcKnG7f/dLs7LUadweHYr/NBq4JAKawCTEgdTRYpW
qK4coLkXjY4NrEBB0a2qNK6iIOXF8Erpd5CMU+vuaeUYb746gwiq5ZiuVJRxYXTIt0iVbOYa1KHa
Im98JVII8NV7dkXKoQ28sewrK1vF6PbF8wcEFXFDI0GwQWSQ1IlgPPo/U5oKFknNPkF68i0i52kL
bpck+Vl63/Nquq6HxV1QwDL5wtZUxrkP97Qek8orHtxiIh/HnbdMzl9SiSYE2lWCJXvRlMMrT3J9
OOcIdgB/wvhx4Nv17dpEIggG9u9E3hltBOwQrai468+GL2Yf6aS1Ibc2XMgW8kxMxF6u3hklF+XA
9po1EgN9YDCBwtDn2yRrQa1I3edE9T71/doLpRH/8DUTd6F21NIelG1+nzQA94VJghbrDjP+/keR
KkLUSJ1wAPLVjPe/Wpfsz5CiAJSFPYW4ai2vZf14eXi8Ml6+cGEO2qUzVNJdMzNF8+qM8JnZh5kB
gGhuOSoLlOKH9kRegG4qqNw3YD9uOfjZWCfYupRF3UbHZ5Sw1Mq3u3LbqWW6Nl8B1tcAjOXPw8yC
VaBoJiawBB1Q3c65g/aF94eH8wLKmgmP0Q5D+Nup+2tRXhpFsIlr6/WZr//uW0V3MhKT0DsqmKh8
bY2RuNf2JU8Eznw+XBsQI9qebiIsobJL7ZJUh1NY9FcgGtLN/ksgEYVpXOuIF36ZrhCWzluWMjBt
UZoTSSOkJkW7ivVAZwfAopt7IfilL9fHsb4y8f1hVwmlaiLw1XAAj42CFYf5Ss45pifLXtAqmwMP
yIuZ6G19qq11pbGiQBoEDI+8jqc+OjPBbR5IWAEG1/nsIpMuGtNzIDrrRyZSV4o+ndpPPxtB4AE5
a4dVkp8xIvDXltwBpanTiJAAJ9MovxolB4yAwsUY1LZ5BNpe5OIh7FKuPxyObsIIhfv6ZHhkntj6
X/V9t2HV/DMzcSmS8Cwwp10zhvLZWvOfOX3AQntjq0IlsXPVmCa7a52u/TNJu/kPXH5VTn2x9Ndc
Pi41YHLz6mjeCYp2bmTsz7c3Ik12Ti3QdLA3jGWKGZa9QrmqTG8AQDfQZdCedFVsl20lvfdL5YiP
FDGyQoQ+BRhCYzonAp1mbO8Vxl63qu9bZm6S7ilWfiPdPDVEUtSTMcG20Fam4QcaGADjTkC0gjtx
BuBA7g3YPKsOgi8U7sMsMCq2fjz5z99tLYhMQvVuOHWuv1u8QK8OTcnjV9HksyvVMlvN3FtD0LBK
ByUi4b373z7uvBEnKfB79lCzsetmjaXqnUqwnIhYN1Mb+Tzg9I2On6Fj4CyIpzIns+qc+6wLQjFh
gWPm9dMpl2I5rjRL1QWgxItb8s9nzd8zKpkfeqRsCZhr9aVaSEW0vCKDJEU7sYlEYfhjzEVdOgJi
pIPdEcmsRUTWW8I0I+8qMEuZvAfq2k/NBu4edmDGSk/wIj8s9ywu7Hxb8iKK6p16bO7q5CDdMzWJ
4nGedFSM9p2igy+H5HGBvOPME6sau/xSO99FsRYCyBt1aiHhI9UT91t6NAx8J8Tc1p68VCPamtXz
zppZzjASR4tDB/ZKlUqFc6KH5XJC/39oax8A7YoLwze+qTVPs1NOyhURFVFaJcnwarfdPDoC/nXQ
NGQanagEaBkLCD3dlnG0/5Py6ZGmYLAxs/nOX0KswKMaArIQGeD9/eLyIygKwYss0lb5Knw/NPE0
MeOywonttxIHIDVIEonHUqQXvQAJTNkIR2SyQTx0MzstM04p2FjydAbYDE+kR/981yIHGg970kXy
5ut4kLkBSyP2JCqWP+uLZMsYcIHIk291UUzUrcTRn+rVdwTobXtCsro6QN58hpkD/5ofn+cj3BNK
9GV+oJYR/pVwYwSxPFnsf9tTB8OLkutolQnVjPIG2Wst3W50HlemQrDYJ8Wv4EIWhRWu6jZ1Ahqc
v42Sy4i8qStzO+KA8RoPoGH1RlRc6BiGqk5kf0dX3G6rs6japYaSxc+0afLVDU9fgHkOf+yfOT0F
o3AP0tgOI7DctaVrMUXth7WejS5Wl665KElfwhwUB72q9Mx5QYN+4QzX13uGAGpcpaBzm4lqZDcP
+BwCk0mYVMkTafasoq96/BU3bq9hKFmxdQPtHymPOiYH0KcZWz8uxn37g8myR2RyDsnEFetMBD4F
9wSp6VbvU5RyUbdvBOGPm4nsBiNsUv1REkyQZ89Ce+efZbp7XvgspTzpTy/DaX0wv8UNRQMrxD/t
m16pJE9BJusISzqMNjmDHTtT0bMUJXOx4clYnKKgf2M8UW2LvsOqAMBad/cb7RbLtMheCHQFwqRZ
CmsYpLG6TxumMZMeNNxrr3noEy9xkSTu2WcgRrh2+rDvoXsjxMUrV1s9N402rTx2z11ViJGNfz/S
OAxl7ZrmIxPqPrMlSYGRlGT2902BvEDHgjsXHTFDPx5RHa7CSCVJKZQtp2yH7MtBUtVjAJMewjMG
Dkc/nljr8RB7OSz5EKCIeQ0/u09CB6eXsF9jFqkXVp4YRurzGrPOFNbo814RqTKV4LC3e1vFPLud
aQCT8Ya8iGf8OeFu4Bi5w3zQB0/gNvetYqIFVAmA3NEKheqUCjLWB5ew+o78u0rgL01WdwtAsCiE
Cfhd8NnqKhgGkNR+Z3Kfoo6H4QjpPLlXqKhgbv2NUDBl8b9v5PTg8stCltD7IZFclVB9tJ3kLXG7
qTDobHZmoVir/4v0m335RDd11nFQD7ahaqeCPALeJPlcX/TQxmD7h/prdA1xdNvffTxOwC1WnfE0
vGDPdNcjDNdpx5jCrFjtl/LMqv7PDs1jZbuVumoVA2ikLa/CgJCG/dl5cxfYteTFzvsH1iQm9BIv
tWHk5Le7hjqgrp72/Kj2+7bHW+aVMg27XDZZudk6atwVDVXp1C7i+iTJt8sddCyaX+gOcV9e5fkN
swuzvQFiGMVq1aDbMnaTcrKqLagLdcp0kdo0zZAlTBD7lvx/bV4qsDSya/0k8+M3Su1qjitaBnb0
SBCq6zvPVRgyfXkycbg7SfFGvZc3w5q4QyWh7BsTs12qPJRuEd2UeCTwXo0Qxio524ckzLMk6Iuo
BJVJ/azlSTL9/GY9gKcw0Ibc2M0Wx/FMyh2KuBVOf1AJoQ3Oex3myjLYh7Z8UU1VyBc11LvUFWo9
b1MQyspu/xiFKJfLRGpfYD5UurE7+V+t/AL6+i4KathS7gamUmj1O/CXRsNGu5u2QhzHA7kRnrDB
W01N3GuOr6g6HJWEMyS3BXof3q0nKYIFCK9Enfcjh3/6iJXpG7pbyZ75CckeQNVDNzFMGiZMSXyz
Q4GrYvzWRmAyMIs0taEw1OUc0OUzHPDddlv4slDCzLVygi8hlnc3gZmq0RYQrRkpoK3lP16Eg8PL
snWBInOhZuNiuETHqMzKa8mNXdS2RogcXLgLGodmDb8kmzOMiPeknmKTjtE8SCNQrJ/c7JddOyXN
0mkbgyFNmzIj+OewFV+yoroyf2WhOZ9igAvCJSKjoKG9DeG+LmJ3pIOfq32sDRWkVTZXOCgncJCs
91kKXowoes4X+mUUIsgyYqLGTTEfVFA3zmUrUXNaxWzZdoo/2MX54piNEr2Xbofvhz2b/eCChtNr
xi+tzViVIZMCvVsUsx4FIuP8MJ4ozN67RovREdL2GJLigjtlcY172EyM2rr/XVbOIpIbZBuFnil2
hBHHA8BPbrjdElhgFsHsfzvHmCpZH3kXWVuOBSzZd2uPknq9zKA3o2e4nlS2QBCRSNcKYUfVRZg8
AAyUgLvwKJGXKnfi94uDylU1M2pJQd8N76hCgBQOd/0VoAouoTFp8OayFeChteWLPyMcJf2jykp4
X2w8Jf/VRtSlroyj88u8rEPkMEvRxi77numWKaqxA2yQZcJvp2RqHTFNymccILqy8MqWDkhgoU2I
MVWy3fVOwlBShnMj0+Yz9tsEJHg+bPy2YZmd0CPSalGRHRF3EKZOnwm61WKrVHTQQnKGK7lNKzi8
N8w8oBrIMlmHTqEB10X8Mz5Y82+ZsbdAuePrhDkRDmPAFg29Dj7utaNiqaWfWmKt0Y9XErKjOJnu
jrYvACYQ5wySm6pp96e4HH040AbknGgMJ1gK8Mlkm/Y0s1lfxNau42QG+ydqrPumzhfWuRz1g9FC
WFf/9jPsYMlSBzh5j9+hMB3Y3FeE0w8qhX+D+M310I7NAhJBXeBTHSeJYb3sUqN8/2JzpksaA7qc
RSag9y3ZT2t9FyPNfjYinQtTZvUvjs3ZGTthYGs4k5hMxPWHMmDj6vOtqwdJm7oK8lTbPJdhoSAa
+4fJ3GZHjeEq3ijckax1DeFgX7JbjmWSE4mAL/AqZsFkF1sWLEJk3vyi82BbWfypTJ0aQhIi3qHx
3f73gcazb8OfZlkMQt03eRL1u07i6q3zO3zvQDcuTcJX9GuW+Yctp75pjS/dyL+dEl0/n8Tyuj9v
7zpGQFstM7qjBrIkclZ+lpu+9yrjab+vi09M3Uh53v9DzRDYDTRmmr9gDDm8GJZkjQTZWpazta1B
nHp4Tm8p1wj8SklGd/5qROYRXUnaFIzQDUsEyOlpQ292ia+E4F/BrdWbUK8MRGdA1ii31fnF9/vu
57oVNA295Qe6tyjCmKPwsXyde2gPH+cSfCCACvNDP7A2xbkL0T63dRGir+Z+7/KT++1f5KGWVFbF
CYO1PRTsD6nheka299Mu4JSalY1BP5uTtGrrVlmNd3EZ195tShCGqUFJPfzkPv63RaqdLQ6JH8iF
WtdDJHlLgGBO1MTG0cocnEu78rRRfzdf4fIqOMx746rbCeDLyyetA8CQbrANBtMYWvl3bTqbIKha
eJfwBVI6tQkAyheLDHHF02AODVqYB3hWQgZSxPXjjNVBPhDtInznMN7pfjBA2yRnl9n/zw2RHgzp
CQYzt/AyNtQbSSzsOv1BKvLZkdpIg8MQtojwV8EiFRH76djdsyonxCRlSf+A0JpptPCX1CJe9bT4
aMuO4g9d9ju2/Lw3OjzaUOcwVX2Wkhe8w0L0VqtTA4bEw23PQ3oy4RBPFefrzUUcY/NcKnVR5usT
Di1Lp7TAWhPbBlGr0pqhuRfQ1lZTR/K2jtr3lMyGf4igCeLt+5EYo00xq+BMDa51ZmX+BElPADYl
5fIpFhovwMGawJTY4/nGpE+yDi7nBBj1J38S2Y34PFvdYJ3KOqxYOwE2lxWWu8KXt/dOYq13wBPe
tQbsvaDLWYSeJABMLXx2BqLW+TdGwbMn2duU7QCFPOKgBnavH8XsDiB95Cu+rc8h3IpY1kQc2JHs
pLAfu91HQRlHZveKsIoXtpeb/1k9bWC8f3FL72RPEJMZ1bY4hUXAFGIKhuCfTl2fsnEjf42bB81v
otLWJ3ENZo37QxBPtmWAMDfj2mTtd1hE8qyaWvkh8B3NOA4TthnoU6uboZ+oaHliTQERqygx6SkC
MAb8O6LRMqBSd8JkU0lum6h0ne24PxmiALu7FHl92fftdgrOJ4M2MTvyOOBF6g8zkW89whrGPq/P
Q5EqdLLz/e4Qv6FhCgyr5BzWBjHE9lnY7bfPw7Qf8JkATlbKlxR60rUWKYB8FsAHJ9eE2841docT
AVXoRlWnnOb6clboSRTJSQd+Du0Q6HKJ/79b4j+zfyM/EPQ6UwkOOOezhSSWOKlFcYKiJTppuaRz
8/QPT2Q918RMpGOG06ptlJozNJbb64fR2X4DBmlISd8MJnQk2+KRy9PhAvikqDLvN8SBjSh7BAae
dRoIzsGTCmsjcKPl2mxhv76L/TkRNctRJh9MPGyZ5H8T+K8RQJ3U1KyF2xFby3IHbGA6kALfL0V4
LwyfnWkr/CR+IGs+TvjlGq8VLef6ewlvGBb5te/EaJ4jagf9f8TB763eWtYDUD9DjWWZrIewdu25
9oJS25vxOcXK9yen14V1PYEH7rPISisTEtf9JZGHzqjTPXCnDeBAOGbyLI8U5aNQ+/k+Rk4VKjgv
eAPLrfT7gORpvGzxI9vq2gnfNhXB4pPndavRF/rMlIX34pg8D7zJadS/GKrrMuRsoZGxpkfciaYo
cqyNE2xwdyg5SVrNQGZGONbJs2NJRnE7ALvPE5mDVxiaYZXrjveY+7mcQ8hIG9ZNHFFIrn6SRgJ6
HFx8DQV1vjGVNhfhuSc2A4rsocnaNFvRmy8l2epZGMYptrj2DMq+9yWRc++e/SZM9jz6KFF+6KC4
1znSftK8nOEgNI7acwttHY93Xkh3UFVIZ/WNNvWrZQvIplmPazXn+CqNh6e6tiaxcx0bN0+RQTb8
lLFsPmbmX4fqgLR/rwtU0R7eTjwaCA2iYpLGeHabTUDxx/K+u/ocZStKbVeNVi6OQnqEwNbguEDs
L1R9FlSwXgdJRzCPSplzyWgdG4e0NTt0ZkzilKlDDytO326D4M8nqKItynFkP8lj4igKb74PG0xD
OVONvxIRySu94Jgh09IzpQWDOsYB4EbMZKC6Hu00JzzQrqvMqz6ZLz2B6C5KClr4oOtImiazIXEO
UijZ/DcpEiYP7g7S+iDB8b/gDQ/DTcLDunuAEAAhtidpvw4mqK0EPZuEqhfaZsG4c+qD3zikMYVx
lNIisaUvIlsfnwaRknrRwgZSl6TBVRNVa8ZUpDwGdQC66ZYuPV61W5/FGoGhIdHnzzVZ8Czj7PQg
avQ2/z1LbmbonN5qi9LY7jSiDArE7H0/X/JX81qpTm58QofyA30MgM2Jtvdsnkv6guOd07Ebh+y1
ucDI18qNdoODiOlmuyzIUN1yLcKt8iVGHtEy+zC+mplmjeNPWIENmPywhnUO4l+jFW5cwNFC8ntA
MPJT1lIgaDVn/qv3mp+9CoLc115KO8sokcqml80JzB1dZHmZdp/HjLZKOja9hLvQ//jUqxWjC6eg
XlOP5Vm14IugitnhHKt5hqy2jdkFI1SKLiJci8SFiIqoc55nrOTaDPaHhM9Kld3lHjfcqnaREjPE
6xm9+X+Kls8G262WCJbSgXKWhjcWc3DJGQPNoomeygv/RKHjKSukASFNCtURGMRihTnlRARKqU3a
5/p/Tuzo2ER7fJmjQGv434ktjvVKqe3LdmyAqdAUyZTK2JqKTykQ0dofPim3EFyLim2RfS7re0yP
eyLJAhoFNBb9SMBTdocCUJaUWZqcTc3iZXOLMoSv6lOJQ1KsiSUDdp7RvsIZjBHpjJfrSSkU7T6+
8R0ikteqsJfguuOo+zbhUTQ8pacOgEcYN+H9ONgHmfwziq23mv+hz02O2tA5wVAhB2XCTcN+TaVA
cLX/Y05j9lLtHWfiMyznq2vNVnLczgvR74+rpMu062AyxZ3ksxPEraWnBncPxhzkBRYIOQi/UXmo
OA64L8HqKNMPQ0sLIwgOFf0dOiLy7NPfiuwkKHs0GtCP1c9I0ku+P1JYUJvAV8yWwK/DG9ZhiYeh
u2uSBqP6C1/SE+xSN/eNgg1w6oplJ7KOCNOdH29U3YVpt1Eao43abqlZJFjEfYYXNPkPtFUleyq/
/VnBZAPo3cpIOvhjEEMmFjzBmhK0pZlGtvAg1PB8f6oJ+TCfch3n3Biqr1/Xa+CglujVG/WnKU/3
Vor4pohN4QRHpLNx8k8yxu+MPTaF9hU7uB7wXFW0nakpb6Rs9rlUivOm/X4VPPe+zulb8fjWFQSD
90v9r5pav3Z0EvWYb1Z74FxcpXqCk5ptzCcp8x2LchNxP2mA3Z80MCA5mFaR8M5S4OCg+mBhcpo/
CpzOLP+C4ns402PBgd8llY1Vx8Naf2vIdDrbU7FgeJA7Uhjoj7ddlDQ+nTYFcqCxMisbxVWFSuLo
tKCVNQGd42Uwa/zfunWSne+rJ8l8XHGg+rdf+mgH7GlPNxj9RGMeOVieJR92ujWNYe0T+cXRwy82
Qt0d2dM2uK02pXMYU7vECYm4rPnTxmTmyLpBYtYm3+xo/nOUK3gxwK90axNRayCWyPhPOqBT70uE
SD/tOUr4ec/2wFF5q1f09G3ULa/3nFnuWtdAnvgfWUfmBAWXnFx3moWakrr93IIXZUDShrmtWvET
diGMzBk8QPmuLiHaPxN/9oDGv9FSflGYS4/AqBwUIldZxxqGJruaaQj4AovpmVApm4NQoaKxlMYV
MJr20GJW7aXXiGXRYwfH8em1NZkv+/glDOgfervnH5DS/9ESdP0wKV7LzzB81lrESqOp61fuYOkJ
CpSkEFcWgOxOgq49IOsK0JmIUkoja0eiWPA8x8K+TIQ3pFoKF5x9vNO0EnRoRp7TsrwNrvuAAjmf
j4tKClHIQPc95tsaoELViadG31cUmF0eLQddl6Bh151nflxuc4fPVsD/niibDAz9Z6O2iP5Nmuag
ZO9oI08MVqAA0Etk6+XE8gK32hTh71chzjgBjow3VeLzdFoWBsHum2jliI0jw/ODi0DvrvVVMx1a
iGn2BOcr1jprcsg4LuplzxZokxa32/4Xr2fXitA1+FBI6hymEM/WeVcIMg6U0Who13TzIQSxRcl0
yogXQ7zIXT9NhIwS45gM7rGqsLTghYdo0sSj+VhCOcVtTexAL12OV8urwaab6g5E+FZ5pfxCi5pp
IJSKFc9Dew6RqHtSaEuLUVT3pVq8+qDLvliM26MiS3q0s4Fzh0vpz2SPvl9zDHXyIznDBG6vUZM/
6JnQox8h4TcrFcFzI6YnP+8rXHmoGK+BTPTNvlPJHewhYhBJdqtUVBy9aVYeePBHH6pptqv8JSvT
+bG/qGJ5jCNzKp+gJx14qWOrVHWjK8OD1cVa46YcOyf93919toC8eocpDHtGgTDj8PT/yRVPuKYH
G0XVvTQ3+nuAoM0ewdpEzhOOCVFK9ND0OWDudmedYWOxZJvgjiCFABCZgCYGxGog5rp95W7xbW1p
cImly62bRImN/L8xWSRWod6ntSyJp1sHpxy3J95plHMNV6Aq0ztSfW3Kw2JQPc6+fvjZBiJFoJZQ
K8Usea+i1ZI2gD1ModG1oyQaOu7+aoDnn26SxygsGVibtRvSdeF4CoON6jauyYMxlPrkKdITk5yd
Vm5k6r4r8wVSGqxLGf8CJqzHLZ7M+OElWdmARshi0EQLyyNNRtyulFljKkEohdcqRh6UbJjqlcMk
f7aUJQCsQcAQivWShK443yGb6L5G0EA/Z1eoSkW9myrspzcOVbmlIvW2FfEP6dWhRkSZY8X6Y1kA
wokr+UlreqqQEf2teyzGEmOXML0Vuger3ElPaT+GWnfp7PEFpEEfJQ980CjzCwPLh0Jq2hq32CfS
wTj7KLyoDZKFTL79wF9dKHApJvereiYBYNqA4ljEyPZR5YgFEAo8fOw4riITmyMpUCzfMHHmmMSF
VkrV7I63K6/8ax115GpshyzIG5RxH6qlHOIV/xoWRQK4NtKny6zI0Sjyh3hv/7+sdbLMtJuzsDAZ
QjbMeN82bcDr5lz/COFlaGMhIinRqRwLzg+BHVXe/x4R4ctFa1Fu7ExBGD6HX0PIpkjKvoIg2bDB
InXdyojwHnEVKhUI6hiaDcnSPlOPTV4uY+aSuJ23QpsUN1tPcSdwEH6gRTOdlXwsy5tA4lHH4bQ9
frMm92Gsnjwrx1qGx4hhAZSyZyAJDR6+VAi9u5AYEMmT+7xISyiSxqOcsv5ushUOk2UsgZULlN/C
qVQZvWs8PoV7KzPZmh1IVuKGbM+NBuk/ukY7+wHpC0ELum5/+Pez98c2Lb0EXtrditZ4Mvn3ZBqw
bUazCSwBVGq9EpoQuCGSminnlVgCQcy6o7DG6F0EaEJytfkxRS+EW7+yVGP0nAY2AzB6PLd7yB18
3pM8NhAv6cIsKjq21uEy5/xP5KqHbXipFWUdVUgYEoGLnKp9q/Hxy/n/l9G53svMW09r6HO84glB
sOCqipngn7sELsrQB2qOWCWE/05SRPAFf4eJ5WOGhWXneRshWIvI1CrUCZD6Ys0958dYEo4bq6d+
c8wmtFY9UNDFjmXwPEwuizsrxUXN5RwWtBG4dNWmVfOJBRqZCw+ilRT6HUuCpYnh4c5kbcsz91FR
v3xSLdMEdw57ZvNuSp3eK19k90WAq5991B07I9sErcV3jxhD+DGx0YYvOxhE+hwIalFCFwZ/ZDsI
GSmAm23Vc7RoGmXT713pj7XmIbGeCnOeF6sMyYlCvsvHV7Lcdaqh3DJp+GydOHyzzc6+m1UYvQaM
RHowszy4PcyWAzEQ5vkkyy0RBIabqtQDorb+D6UNbcCVNBcK8Wv9kPZE8ZliEO5Go1dzJ6LLz7Da
j191HpxEE9OCfq/6dhp5NEsH/L5EscdskMF2kCC7pz9tvVublQwAD3p5UGM2hvLJkpOF7BTNfTbF
2APogAzgPJqFeKwxIqbeR87iibLboPBEOJgWjQkXmYiCMHMR1CNLeZmGBL5XTPwmRhSucKWoZqUX
dVvYVS92PxXeOfTw9OBuj6nnEswXpfAo6YFmALkNi3KW2n6YhOD8gnnyuB7G+v7QaCO0IN0TMCPN
vqG3gEXbgbq9cF53Yt70dFPgdqDgLHMUtgcaOiOAtb1xT3C4dVXDPNO7yDycJqTw/Qy3pgsBOu/y
0Cbi7M+VWctgSTmHAqYot2QSjE8295JRsS2ygJRBO6vmTVpww0vsUmOueP0fZgXM2uUrz6FkgtQa
FfcBXVhAabWWbbuUAs9MKaYEH1y+vVMx0cra9WsVxLMkXLGgHpEDl8sq54PekyEkpxD34YxONsbL
aoNQumCr/Fp/XTW+WOLZctEV3rsyHYnzDvIjn1UI4soZRDUpwKC+2dUMa3mjYtcis6PcirySKZ8c
MwH07KrMSeJHNUEeRz7sfv3/M2J8GB62EFpkoZZW+khVg2vMBs3PTJI+2WrPw3WtcPzgQ4i/Nosq
2By/y/kwBs56C5ZOAnElHtHIJGv971Fadpo/hZW1CPTq4SQMwBFMp1O8Gvw86Kp5POS71pxRvEZq
t3sHEbaamDbwGGxzZXp/T1rd97s2e7aAQkvryAHqp5EdGPlLmPZCwYPf0iay+5zTZEziRpPdoaG7
H6rleY6AIpfGjbbxaFnSp2hy2Z8LCEJuFymZsKq499P+e8rNXP44x0QttKIJpetFubnXN0Zs6fZW
3HBsEtYPjttNVANa6mwS43dcZrs8xSHkV5vWW15hgaI7vNl7JsThsjlK57FgPKEwiZ4eKGa8Zboz
usq5gY2B2HvffsU6cK4IqGUf+xe3CGo0/aXiyVXYpgX4NkmZGsDvsJC46g2VFM1+bkiS1pYQJJGu
HpbbUF1CToku4lSo2z3xlXtZ8TJR1ZNcVYYatYkSCjevZ29zgcbhmpJFJViGN+GitULD0GTWPthf
Kf72p0++CkTKt2aapi2iCeWNjgvl0BFlHbVu1jObZ4UpeNSi2Ncaerfj3r4VZqzdlgHcvpeVR4Kc
IOzRRh0k3AnYv+CiN7QwvgSn16nHKbROBDA455zJvO+4Sm+opJg6bOarURmGLxBlfiBe9qCItXfE
go9CZ0RUxUqv1Gic9LVn81wksctlGf+n8/rdF6sB1ZdZ/3Mdrz70ptpczU5zgLJBQIOQJJsaXksX
HPZQb8wcwdWRDz2lgYYEwctQI+rMBYG7wOwK3ZInH+N/pqGyHLeRSFqRpbBvnER3EAUIYvTBpVhw
9a6bdQe1UGQT6fWfqow0OpYBcE3zA6vNf8dYBafZFuoSXACyovfRxXMSks5HGR+3CmiqkwMRJrJz
zjgSLc1R+8ZPN7JwGNhICdmQFMbl2X3IS0QkesFJ2ub3gkztUnRzRxSkUd/bZMt5fzV67T2jedlj
W4U3PPgODWJfjGnJRHmBoUrjCbkKqEquB0rJ4FjoO3FbnbQ7p3bLQxH/FYcQkEDGocsGO0o9J2q6
oWx3amk5hvwHDZuR7yEhYrBVNHkNy3ZoHe8hB7l6zh5ZedNhmCXduVOf2krvxgdmJkfa4+fbqgBZ
I5+n3gGjBTEBH/mB9PnBeHY9bd8kn8R+tjiUNyobmPbGg6ama1ft8FPdFbbuHIfe4pzvan2Ow8mP
c5bKlHxdPZ7KJUesRwdQ5rpKjuuZIFcqK+ebTNr8QOwIqGRrIuIettvM/T+KDW0QXodf+qWpOL2O
m1hIXlnPBIbIypSNhSp6fTJb3T+Qy5FWX7U365NrBe5J+gVr4M8Lfi7YGapHUDrYD7DbE+CKnKi2
RFvs24nyq+CyNKlpGhE+B0gvubscPYmPVNZrgLHXfnXansKbHFVvkNzco3Btphn8KlOCaEeXs8+D
volAWbRy9n3YpMR/Rdp1lwcivSnA4itpNujTcFNVqIYybweVwIq168XxaGh3wI9Ox7SNyNr4ukJB
volurjRSaoednsrf1p91ARHm+2MOBtSrY0XCD47QuBGe6Eb1AFnqIaF1tpiawvlFeFujoEYeX/pZ
DyS8LZbGTbbl26wNJoU/GNVXj6px1xUyRZj9bwkz5bdbpIli9ngBzp+T8Jih/8XZVp9CyLwNFTUA
QE+lN8HzhqqWA0Ab8Zy9XPUUBB0/mfIDJFYrZQ+b+Us/zv1BAmgGPc0VdL7//RIiHKpbtHTqvILE
9TMZy3+BGujv5LmWWCmh3XxE1kosIidNn3jNQK+re9SH84vEtVB7uRCkpsfCG5cehdX7wLBmmyCN
6nVMOSqK9k//XRm5XEBC2lwOFgH0e1hVdb+LORB6jPbZ4p+Q3QNE7qujwrgMwdSU+akvt0foSJ7d
xFpXDu4Sum1Ulnsintz6/+ipUlzQc5sC9iepPuIhWgijumxpMyFkXbLDAeFv6KCXY1NMb0KUeQmj
/GqypH4dS8gL1vkoG6JJhQfrcgkPoQW04zACm/wVyI5id75oM8VsXPAdbgGUqqKMluBzAmB6h/ha
AI5XZh5Z9w6PF/yyd9CE/xNb34m5So4yLpnlE5bri/bAo/B9eg179kZ2c+BXbEFH5yQXsi8/uGNk
kNtQxQJSYIY+iwYTV7M2EvQICMm3UtrDwplJlmw+4/1EOIu+t0FWjKNzMmJiuiSA7rQDjPp2bJ9D
LTkv4FHhCaI5lSelpNAufBn3ddF5fpZxeO8F/jejSM4Whhuh57nYKx0G2Rx4HJs9wI3ispJ32KEV
t0YHLvNE1XbpL9muuikfGUU1XI9vOG4vB4cqxm2xyD+gdxeiv777Lk8soqwqbdFBfY0W5B8enBw3
l5gxyyqgwDgrqW30jVyYnIapuhExId102mzK2gax9tMznvdvwlYDNtSy/j9fyYDs1y3b+HYs/q+F
mEux9onf9POPFUMyKuYkwPXUus5iEX//4X5jDmTzU3uhrfdeTNfzvYFTgXB/osXKmmBJWJ6T6jV8
v1p0swvKo7dQdTL0KDqnonTt0Ky+yxPOlsUoJ0oLM4lHHc5pNbcGM++2VYnxO8Ilz7ffQzeAIaw3
sEq8VJ58HK8+XuoRoyu7gviqsFc9ha3tggvnK/KlypBA6XlYNrjDc/5xWbBoNyPAcjqbUZHrVb2Y
Xqtw0W+StltY3jyeWzNZvk60UQOh9VT1ohFVgd1bXtMC2NryD6VpKG5WYwJH7Uer+TNJ+7dwkvSh
6V4PIjHIC4QLWHlTjkY95qdqJn8cl2631jXCCVYWxXXbCyldcJJVpXfPzn3JNfAJL6/MwWJyiPYn
0277KVk/m5ENB/x4d9aqBw5NEK2xLaBXWXASxFWzdE322zO3vZupClFUusGXHt8FtOUS0D20kDNC
BXXKMs6cTnQsFtkbh5ypzgGQU0Yrz4lvyDJaceo8Yqt7PuKQOCYEkCKdFMStkeGbZI/Z6JZ6dwKf
8O/8ux+rk0CK3qZLS28jZTdkvYlZCDfOtqvZvS0zJQ3hZWz3Yd7+onFlFGaH9DFy7uqx/YbQpWiF
MjUI5NDIiDJ5wBSMxP8v8XqdQdPBF7Jn7ydwktVz91ZNV+pxmCWcEqFJik44ooTnLuAgvWeCokkO
ZfaDjz7e4egQ+CMqRvtbArsuvqDd3XSQ3X9cINp+sCxt2BcGE/g3zIXxTsHOL8PRmc1y50QVp26L
1C5lGL9c2n3gob5OWwVsUGemstP8XYakU6Uqjs3s8VweDmBtJ2ZT/4UUnZg8bgMa3K7lZVt4rKYc
bNBGY6bvHfJJENLigfZhtd2cGAdutYz9BvTZdUf7ZyOlw1wB2N7p54Qqekteghrm9qyrOVQORqFI
8pMgseUMNgc8fQ6R8vYQ/Hx19JUE5DQRjVIWhE6TISJ9eMcmt5BnxYEqDDVlhdba+sP1hKRA6ZXm
Y+7urfqBUDWjBtAknycA1r4Cr9Idp4DCLWX1HmOVidetMaa3n2gXbe1hW9wfSqzMvAwgtJ+sfpHK
1UxfxgmW18Tz8suQeM9l+Bp/FxyRbCFVNwmk/zzhzsJkkjVu0Fo5FPdmtuOW59yEGA5EuUi+BQqm
RFZrII65MNhBZ2JG/IVFuBhTw0n3fk+mau8qkfvzvQM6IkXoYGN5NEsZ3dcZgPOReiLxPFG7xFob
P5KpRt6M2ohB+LBVyaXPnEcf4ZrEIouf/A++K+qW7F3iko8gdFZzqEPuBhKhRs4fWOHqQQWrmx4i
5th4sAR+isChoup9U7L4f+ZUfpqVcaa0YW8WP7AFjQeoUmY0ENK5eFJBgSehMspFudaSGqYCd+xL
4/QbSbnnAfp+CanV6y9KpKK00qcsdYtl9mDU0KLqdTK6xat3QfWE/jV8+bXVphh9kIs73UpSL08f
SCbecxHL2VPDfRkp8xBCZQTF4rGfdos66HtEtjMNepdk7FMXDD7ymckdWZXuqTvLoEqg9PQWD+u+
eGzVdYPCIrinhPrcZpJqfavAkLTSnYUEwotm8012og23yHx5ddifwiIzLYxm3p9VTkUGqEzePp2B
WfGVrBYPHdk+lkWcyRq9SbUGDFZ4Bnb1i9kbzZfk6AQoll7nyuJSZOGjg/7BclOqcKMyXFDt43bD
tFtDDreguV5Bwci71UlaWfH/ikVvn9HGVBJWK5X5mUYAip/R3ADz/JneJN5iE1k1Nq8VP/4vDI5w
8QHW2bcBwYeGjuNOEpwv2iVVOffaCZ7xV8eY88+CWIhaIInwK568nj3ivxo8iRMPq6coLqK8vGGn
X2+IFmlDFB7obW29WvPJtKdICStxU1md9EdwF2/O21Sq3eFaq3eTJQrEBiRVEqb6X7uKTjvlVjVU
CHPfEpp2Uc9E2FhYhHbkU6x4nQeDzETA7jIPxrdtPBocZSHfQcXDfvOEL+iNcuPVgC95EPVJ+XlA
HEF/tf9hQofW3CAZ2IU1tNm4Ob631678Tqi8ilAonBnf5mYsZKNVqY8CRJQTVwjMLKIjFCKTM4u4
s7kLrbV4dNW8QhGjvF7p9ATam8HHXVl04zltpYlzjqTgDmBWrcyqfmQKtsL0EdMA70b7GEgnEtCs
4vpgrAj+embF0tPpGsNDgnEf2bxTJR9CrBxZqgCuZaq/X7ut740JgQrp2qtAKgbD81950rwSjytZ
z5InaPyPNMQayF72AGk2oM/YhnOpHJ+Hz5NwgPeiPJieCYHUE6KzhTYz7iqXQkiieSBHZTbHPFmR
w+D2ad+XM6Icm+7/4f91+3Kat99+/GtBKuOsosXhjRe95Wu42ibKiLLnjCnz4Q+SLYEX2pmfy6Wq
D6pRZOiy8t9TgTarBz00YHLpJT5piD7CxkKFnFcIUkMRyOwUxU2iVXCb2jEuVOANl6JE8zRj27Cm
SdNnicak6t8QGVwVXA+Xq4R2nbhA59T3PIQ6jvGUOrH1qsF7QupaZycoZjhFTwzsPrB5r9AclyDl
iWWITBm8iWnLr1GmD7NQ3HD17qrHJIw/Byl/1uWUBJyWTKTokW4vB/t136UeADLDJj8AD8ziunXo
yBjDmifvJyPbNOkU8Cz98e8V/cBxbDzgGtsAI9XD/yz6XleQpzpcWByC3mLK5+Jb5KwTE5BxJxUq
5QqbCNDPi+DYidcf1LaAXXKC4y1Gb8sNMCfLlL0CvkYNNl4nWYF3NWZWSqvQNT0+0E8s2kfRY/Bo
A2VV70U1sPHj+2CEDsQmNfIOcK0fYO/exL6+z0jzBjcX0jq3JeXincsuOvtezwfCxuSso/2LZBt1
fcy4tuMs3eoq+UjnE8mai2BX7DvtIBrd5FQl9rxLG1KqkR8QT2XlNSarAuSU7s52CzhS+5P5qDXq
4omSYyGBlZLD6iynakKNQc+FSqVLLanVLJoagqJLtYvM+J8OFW/SWPxnLqmNTiP7/KOXg7XBafbW
Cv47stu0HIpeOnFQgN26tTIqklwspHINgmxxefTOX1op0nF6QEckU0N19FrnLsRZSbWgVxS8HEaz
pev4tJAjI4VmrXOs4N0VoSy/2R8S/eIB7aQfgnradLw1XN4kDCXGOY4j+T+V8SthZvDeOkmx8mEn
WLoen5qMB1mfuXGXCRDGhwFtQx9iVjPJkGob4s0OpN+1YoVkWGPs1WPjhYroS2NA0A4kzyLvfLr8
zovCn580ZYBWdNppBcMA320w8aeSMgOYm8bQ1ksnVpNyh7WZpzYBnSIJkBT+pukFI6CW+OrNejZg
2lu4vopbJ3RVC5rfaRdwxaupf88mu7LT3aslDP5TMxvaqCBjDAT6clQLSU6YvHb5QVhhhCELscRT
pn6Gl+01uNP9P06RzCl+9cbEW9wcK7WqCqIl79jIzGf6MeRjUzwNFNE7xBx1PoPM8+wTNd7bA584
OrmuwB70SfNNuhlsOCUfvJZr2p0YUX8kQjCEs778L452RPGqWRcTg7Og4bjsFxvBEsUe/RTM1itm
F9evtgZ+Ms9sUkBcwY+l3WDgBP/QWlHdzc+R7O6+kV6NWzqzsdHTlq1tMhQI0eB2flKDOOoz9HHf
VjqIOPPDDR18sBe9zQg34wO3v+Idki89551iioSiVLXwLsYRTMQ7iySUGbQfAo2XlGlk4QnM1tDK
Y3X1P7QVcosmSiqT5xGYR2dM/dNHVLsOHxixfRZ/i5+S6asrinpfCjGK1b1DRQYZM36Ubb6Z7C1q
klCHibsfdCwYvVQVu9hMuT75APX0IAMgPHRI55kcAloCHoh/oCAqDSGYZYMoKsQVNXPH2k2SRRJg
j/WJ/7jbvfe2lN4M2tLZ7NfmF+FYqTv3mmRH+4/qSzcReL/bn3Sym819UhvP+iKWltiW9qOhiyO6
dxLQrrpTJWUWYseWpW4YxzAQrU8SxCbZJWhP8XUI9GgfyGqHtMksQjH1EJ6TNL7yus2wj7LJ8HIP
8Q5KVJpY8bY+me5exdC6sWf7Yj9POys+i2PTnKRuC1Cm1DpqkzbtY/pla/vBkXF0sRl3ibp+TkHV
dBFr9j45GwVqm6IewLnkTWSnK2YytJk2UfjcpRoPt0MQlqHfNkPM2snwJMHKZ7wCFX0nztOdxvx/
bZyKqhwZVUWm+lrPjXMal0Z9BWOESrrjt3QgqsPbu3DzIgDIqmxj/MGuqSbTI54OURATPX1GDyms
ONWmbvWD9+fbMecPYCTVUkqPVUMgKI25GA81PGEOtu2rhhX2PDGAtUmDM0ccPLbRj4IcHv/08WtJ
whP8p//0utomZ4IzVg3SmrJAU9iVh+fdtKc8NYWVoYSwH4brJl9CLCcGymtHqxiNl5tNwHaqAJ3Y
BcaPUWDV8VHGSVdEgE4193HYd9EdCxB3b+mZfYviqjNZ7oP4ww/6QwXWm3j3ztM+TaN20nKP9TZw
v5SpL/ZE3tAMTUBHRtrYOnDTjvRJv17JfPo89fuco7S4pUP6iTzLtA7Fej3lOPJs45rRRxfwVDLJ
qmQVZQySLPwJmyF6AYewY9Tci6QeP1WnoNDm8qrCHCiHT+zcLN9oePJVijSGgX9YmoN4c4D3JbAy
ELOHaYVWiUeTdSW/USgrzWkozfrQ4Ef8FSdqH3rT7wFjmcGFAwDUoAfYdpoLkQMwZ/6VH79Bj5hP
3jX3qmOCfgdpaBQjmccnj0FK+jYQyqVptQpAQlgBh/J5+gxy9YK188lmPjR//Qe8972yecyly+hP
qlcBE7Ymy2idPmENgta5wo8KgcoZtX1VdOh8pnSND2yU11JQgMlDGpi/uJsIiWzSLAM6khUcKZ9J
J55XLYW4+/LKXefK3gMwkkFo6toHCz2/icmJfxpDQLllW1DkZkakrgX5cbsmMWF5pazVxRHn6DTG
orPlxhekZBqCprWKl2i8ltFEzc9vCtQ4KUaRI1iI1lCQ0UYw7WT18L9/qx/8p1Cm9ou6ILyDQGkZ
uPCfy942bamQk4y/5kTP9tve51DnQzbh1ArSMnmoYpr3hALGZx9FWMyNpOQsIJfCbRc8DcR5TwYm
FB4spBAhQM1Z4j+nu0obEr7xCeQADk2xcuwkpHi4ubhebL9Az3M7RZBzNWu3P2LCPpNNpwEg+hyD
ETBIZH+xHjpooAY2sAH1LWBGppOntBbGiP961TUIpZwX2Li4yXUEro4OJnZOKV/P+JEhU3HOpPib
ZgkfSdSuvI09v5yxj+DbyfDEbcgEOygfvZgaSF1lhH5lQGDNOX1m8bTXmcc8Fb4gha+uvET7xET4
fDMtiAdtW9igmO3QZQA19F22DRYLNAKx9K97IwZEFB55XmNBvfRRLY6UDJuFhHXNex4oFfE9uTNJ
CY8F5Df0dxAywUrkg2ZVBBwhx8YNUVHChfc4SxutgGlj1Ku2fq9dwHiibX6W9x6I9UsZ1RAr9l0W
NDG5k9AlFq0rfUasorLusRXgoE4Erzm5ELiDs1N0Ht1lBcgk/lKF2fCuy4Svy7XTnWgbTUHpmHW9
DZuy0PTEe3OOpR9zAQZQqhdiQ1dzS6xerSbu+egAHv/FuJdwvGB5/+s3tfVrGx0RGx7ld/nO6KhN
EiKsSQG0bs7gOkk3o1qSZuO0aDqUffjq5fNyanCLAVa64eDQP3ewDym5P3FBoEEi/90oYjRNFeqg
mpDW7o/PDtDj8MLJdWvJsNnlAOqOV1QNqtJq1OPf3gs53ytLcGzW5OuhUaLCbJanQclDlkKhfqYu
rlYzlhJ8TNJrQv0xgE38yMCI17l8lrU8saSeeZ7QYfGeEAq/X8MbC2VQuevZGsqpr7MK+CGoH8xV
wVY75smm2U+DblPTgyj46o/qRRf26rsOed0PV3d12io3g1CUojcOmDMwjhNWZXKw8R/Hqjqq2EZi
up53/WONdWxOFxbfhfn8GjkZEFWI4wag+uKFj51QWqCkjFCMyQrv0yAsiFZwjCQksTluKJ10eN82
k/UCDIqjS6RaNrgo8wRSyARJq2msKaWPoUV6/Wd2T3WfJMf19Yl0aJf3sLaHFVi8OR0HpLmFc3Nt
woLZzKEiyri84Kyb7TZN2rsMi3Z7e9Ys/yd4wafrepjCbxuxrj7yRDroyx/h8ijn1Fc0VHePiLbb
IoIQLWQWvDeCq8l4Mw4sB9Fx2uRARUCCHpK2I2BI3GRpDZNF9+IX9rV/0/zZ2vmEdMJ0xHWJ8rGi
9MeWCtQZ8W0Jz/JU1L4o5atwfE5RJnCTlBOK0ZrA4l01gx6qlpusguNYGeXpwjthTkkMaBGdtC+K
6rOPBCjVlxTJQOYag8MRZf3Uk5rCfAipVoc1ehVt3DKRtP849HwcCePYT2ml5deMt/OBPT2G57xp
d8IYwkD08DDgxQzeUY49BZco3SK5okIf3K9u/x2rQfcSGYt976iXJarZqyms4WLi9BEE9euYdV99
PX7+ckBlzy7lQ5Pj89wapkUmDsZsm0mNQG8UGC0isACOYajQBqClop+LVYuNzAniBkJDSN7JXxwt
P9wgeIfPMVw4+8r6dm3Ngzq2de5fMn4LnDOidIK27kyoBBhXdUPwSPW2WqkW5VVuhrfqzFmi/Xe7
w6BPzzHGMw4+i71T+X4SaVrARq6Gvg2WeeQt6hdsHjALPSaESTrGDjEUsnk/oLKjMz02uyVxi9qF
FrA9yikvdaL6D6GoffgZJGiLdGrGrLYf7Pjf0Kz8sM+Y8zfoQprqc1zeFcAbkqDzTybOz+7blIAF
/kl5jT5ZTEFUzkmCLhKQLlq1RFzEI+8SVMm5ReGuW1dRGYQKSrp8kTR5Y/U9a2tMDA3ylf98de8z
tpSzMXpMdbosA3H9EAzv1K+8TlqXveTxi6aM89G45BXjXrYbavuqGJWZ/8PGoTFBErzgQ8OA70GO
1CAkeiBPt1wcBi47ZUA77PtE9emyVJBhwQUbwyuk6JGuNLKEY/IMLimfhsVq8fXz5lTUwF+ZGUQs
KGPlOHKuQnvsn2Wps/elYDjNiD5466JZRqX5yQoWNbauAxiEsPL345fq6ydpCG5/nZd4KBABLc4D
94YFo6xqO3B8orfwjdaZmB3VoDthDckSa95JYEkvJHN01+dgCrF50pla3uOBqa6RaWgSzanZ1dIZ
9c4Fq/T++6l2u5uA5rQ9kF04bInLmRnpRgp5cBqtzAzTiuYM8XdhH+fU1u82U8fBK+1goYwxwwGw
1DGoAKw+kFnzheUb3ZP39pZE5F+bHa7X5wPQlwtMeBEMQVfdKxJGsLxDGLNkiGJY7nQ/Js5HFBOx
ZL5cis5izJovR1j4yrflfdDURBhdL3Cq6tpBxmjd2RJyUh2jyXQEWOmvZjP5wp6jqQMBv0Hzd2ba
RD6QqY/U2w7GGvrC3RHjmVssvAMP1lBKgBeJLUaChXNqq8blV9Cak3kgw7B5Hy0Gp5wbVdT1Jc2P
kkZYhHvhbS8VLcNSF43CDoMIlJhI3gzv15Q50NBCXPiJtL2ldbhPevZ8akbbcaKvSPks/Lnwg3Py
ltgRhp0Y2nogRSDDULMdNuaFTfxp+I6jADGaN2bJPFY5x2gEWsdTRfCjQnO2rpKjPmIqdvhXj3SF
DA1uOVXeN1xedDRoK1gAtznmJV/Hhn/ZpgvTyQiwJb8QjbH+Opp9AcwtwOcF9zOreS0m4GKw4ubd
N1UPJpIXh4jSqpkVKbkIQcWJy9XO5EWqVnW17q5Yfw3Ow06HCCoYbPq/zW9uxkK9BLolPe2Wzy69
ySqMNQR9ptO1N2tQ5G6oBdYTz/vbIi0RowRCN2BmHshqfsjZwN1SvlifNOOTu28kBDxo2xUJj/sd
wEt/IzEJEIh/hKvjHeM8AiKe9yCeZ3cPhbrYu0vbWCM+UFy2k/AqqL0rI8v8Xiwbbl6Mr95kr8U1
THWBrIdNQT7l8vd/2qVHEvl4ucc9nvKvls9VHWI0I4zyguslYcpPsFswvT+FaxstkygGbK9oUqO4
oOfj2dxPzzioAlr7a6P4nwr3EEkkKXII4A7EJYBsOG2awb09mUIr5Z6eAyzwiqNAsiKeAxzPtNn2
KXg6I3GoxcdDxBn+eSj54b1xt/Nuw2Q5pFJhSl4Msaiyvxp1TnOTxTjgj5csk4j+0g8+PQYUUqch
oH0QI4eUBe9v527wfcaieBGd6FmYESNoLNum7DPPu8mTBPfXkyf9ioHycDdB7OOF3KTCIh0/GXXz
4ima3UaRKrrXHgmf9W5YElTZqvhLPZF2dCelomkHCyX8G6oPmNg3hOesP4pt7WsByOYEmKkQuJ7c
TKY14h0p3qTKdXHxdnfU1LT9k0itEYDZ8P71BRlrgW+SrXh5IDXCLG4uBC1iCJarS41+XUW4wzso
hW/X3+WkCNDShgka6/TJReh9PrpFjiDoL/gh3gZAwYMJeDGg/Ur+rv0Z4V0Dg3p2qPqsWnINAGWG
IJ99RrSK2vUUefjmNHBnQUVeRwU66DRW3t2b6Tzrmd3Fv/PiSwAnyf4FENSQaWM63XRmxhvlKP1q
39cWpL1d00BdsyOZ/xJyUqxX9ZKBNdHxVoky1WI06NnzpTzMoPsRobbgYlRRN2q7DIJngQofdwQm
PLFwjgzBKG3ra2NAsavo0Te7mGxLb1Mn13IIul5d5elvt7vbYVf6EhqHi8v4ewUOTWVIHsxfEyQC
1Xykv+9vuuYwOTJjZFhJGN0e8hnw01fpyDhteru+kuhqwZILitX3jS48N9ebIGB+Fd6XRHOe6Hhr
Q9EEOxunnfYsaBYTNlbFryOSG1TLihIXYMvMqenY6c1n+O1UvXig6cK5mENLBlYP98WXa6hN5A5r
jHUnr6wvwbwyWu8HFDWZYhV/uQEbG+vN9UrYeiYdzhRO9eGWlAEkzoQKVO9ijI7kjeMlzDHpox9n
kHAKF+Pv5z9Vm7NVdHOTTvZVc/mxdy5K9cNBfbZJ07K3iP1Wz6hwJagpYuXaHnfTIIn2gHU2kWdB
vgNCwbFVkMSVp+4Rm77g3kmwRStZQT7R/ywoCJYhe7zZymkeapzUZzpua3EPCJt15RYB0umTACzN
cyCRyYfWcqHFx4YcFEhnHberJCIMyfoT2cVFcuhVfrZRh0WT67PN3h0p9LZqUYQ1kdN4hZY/4OF0
E4/dvbfOX7+UHx+h79oq6ZxM3Pqyxz5uEblQeLEeodEbB/YtDUBgGQ1Tjb4atnUjON+yxiq172BS
i0jKq4ROG9+a1xlZJ5I2JJrNt5EvANHhW2rZxDtgELrztujVs/wRjDRgfzQ0Ilh3vNlcEmrcE6IK
ye/V7uOUPy4u6yh0nIDRBpT/SGnQ45IcQlzkAfvDf8GphcVjCROaLe280gldTTgX7NQiUlCG04mC
dZAg1eCG202ubZv31XJP4tXGD9gGzUp03Rb/0GWjIyq5q1lkuC90o4CoJ6V7CCJMKAmKNSHqV/mU
dPS5d3IKzn0lxp2HwdB4H7oQJSKfGEaF5PyWbX4OrS+W8Pof6mu/2NG0Dba0x/9DHxbkSa7GM62r
5//tKIeKIhTLgyQQXQUIQeKAhs8pTsjb5eJgdsc06ttsOiDNICoBbi9WkGXTqjbyGKIfhJ6oX5IH
l/KiWE/X7Bw4/AN8LJEMkt6swm5CoJQ92D4DIO/HG8yrZcBa2LWXD1TTRTEzX0/9VpG9B0UwoD1e
Oqoll/O57YynTqJOm1sYEBng+sV2sVEPq3BMS3c5A+9CQnQMFqspbAhk5RWu0pbugrwzUOo3Rhft
DUrtihlSeYTt+IQGptjM6lrJtUrXfdI19GaqUdEHQLQlBrkX9WVjo5QRPB2N06whboV9folMWrgZ
T45qIDRVjJS1IDvCUh7Ruxf3V7tdH5bGbvHHRh6mJqdagNXA6YBYkCe10zuhyrvVcj5PsD2sFHz3
o1JU1LFZyRQpPC3/AQDjTUfw+DBktMVvujGrgX7tXifADU2YCWtPudTXWPr0sZW8mASWt3ABgKtK
Lj5JY5AuusPuVZYJ9QL3+u1YzNSyZQDSj17pIRiH5CFYPg7MwEOhtPtd6SH00BpjNkldYE1jEPJK
qOnRgxTe2hTQEcWFl9BYBTYIGZrj5yIVaeNBGQgXr/aFXC1Vd2vknFNt9bT1VrN020QuDlzB9jPL
OpjKs8E9ZzZ4s7lEQjwHCAYNXEYZy9Fiab7jjTWmfo8P2Hbwmb8TB3fBK+Wlw9UKHKKc2AE/big9
SUN2zpZMENd7WivSIAqi8ZET2aKimci1Vka0b1ji2X9kJZ3UKve/CMhuhvWt7FRccNF02orRUNyc
TjgkvIUD7EM+IlTM33gPLeuAc7Gq0e4eW2+ThbLO26D7+CMkZlNp9BDF/HHyN0kcb4zi/2BlfdTD
TbzoZvpi9NvbAdNlK9yZA9zP2EQ/A06k6xcxk7rVnjfJFJVfWR1xmHgKJMCIo6RVEVUWxl06xcTU
VA5YgNtM49Uv/5WipUNT8ydi4bs4k2UUfFLp4iv5OfbBK912OY03zRbs3+TWDOHMlj+fVQ16g5rv
IBhqrdZpO9eCP1mxZHtpi2KKulCZDpLHwOcsllVwW97Td5O2kXbJjvuYs5sx2TIruOxs4029KrF6
Gz1x4nVrgXwTp1bjx9nEILBuJaOCZspgfaaUjhra/DPwovQBKacielJ5VOg9R6ibETMDYU5NfzP1
SLb3XB/vOkGfibRVaQD2U5DonGYnlrc6x1FC36GMnBTaak/lK3sW+N6GyaRLeSbVPrGeFrsMru4X
amJVlcG9hlXZK+OcU2uYa/cQAndJmCY1SfPCfG9SDY16BbgaPhefegI1v6sJ12YaClGI9Y1R93Nn
kGFKKnMtF4HuJjaK9fqpw67ow56SmJS9HaBMQA/VrPJIK/0nuZj8DytoNArIJ079cj330ni6b5b1
WbH/vTbGTNL+SCwroQGMOkXUv7E4UAaPop16ZFzPYrNiB1UXHpAZkPSODd85nClqKxvFKZos1Y2g
23e2mM7YcVVzzGWQirhHzIZFaHekSJ7ery4JRxQH9rgmgx2jjgT3lAaBdXTm2021eHCvM3u9mIUW
gNkalZc85FYf8Ruqo8cVmHoZuqpCq4JeZaZcqEO6fnD8O5kXoLjfzjKM4EsZxm7i0B2nA6/ELR+w
l6MoCzqOcNMNKyh32NDTzn6ywaysbRr0RG3UsJOAMtVleKjBPWX/AntdDbPK7jzur0QBEzp6CAe1
suuK1qX9Rx6VyRfiFyxbkztnrQNLh5rXGCZRtlSAEP3iT0Mph2+J8nfXfZqVlR2jm42SqO/5fCGf
93pQNZEX/cicJxr7bUBIGCbcXCx9zJptvMHoEq1IAU8CXCPk+jmtBem+nHvjwkC5+vJ5K1J9v2du
NvNl2NoX4FnGs3s4IS3hRVorAqsIizleu83SPctRZnRj4aei+nt1U5480vZdcYJ4wZvE6u36KTu3
1xMa4Xkt4OQRcf+OD7mDuITH3wsHyjTIeHo/UtAkuSn7KJ+vUdkgb4zcFTYoH6U87Jbol+afXE24
cCdZ3xjgH/wSV9wn9DH7gB1X+Il3ZnikqxEyQT6OQPwMeR1zWmEyQ6x9X8+RvMKvIfuxu1GXFp9T
93qQGV1SwpEg5uhgNEQYbTkakIx9VE44grhMtyKYXoF//ghwBI0ay5tZBd0EdTg+5V3T9iiBVpzK
p9/zVeCQhkEXgtblTtLiclQqZKUd16MY1dcLPefRu/Kmtz2oe/Aq1uu5y+S4c/vByDcrzdlEm1Sz
bZWGDZaycju3V4g7WCFlXNiAl8aPDfS8d9PC3Ae7GcGyd/8MxTuie0T5tvq5dj5rXuHt8l/cPvBl
k/fNyUKf/iyRg+jaAYgYBPUqCbJVDAea+0MHVuYVCtN2a+UL3VoUcxH375iv/iLSJY3gg9sEF9tA
c+xj45AmS94CNXJjIwpygJa2qjC9yt8dgZJ+metdARA6FlqR1gtAnzfmKYr8c/exkyimqUpT1N34
Hn+7706JBrS/WcRmB4LIF4YEVMcwuBmDspKLRj+OVlaUjg24b7Ee7Y03fj9DIviW/uo00SeFgPD3
3LLSVlmRVF1RmEdN+UAVw6BfS1UNTOmXtTeV5Rm/n35LlgdTB2c9zeEdKP+5ClD+9pCE6ooAGJK2
NzwIK1UX4yuNXa/C8uyKVjmjEvaweNkxXydNZQmbYTxyhOr/rnMt2tN9q2Zw7BDSTKOchgTHsNN/
ZMPRwUPVQXvfoYjtuEGxxKH7eBK30bm/8FJjLeEkxcjH2E13ELLJT0Hou00RneRnT967tPL8/vcj
QKHTtHrcg2Jf6XpYYSQpQ5pns/oePgQ9rF4kKPU3jfd1jFRDBX2N6JVRDwm1inZ+lf28Ka4SOKaO
qIb2Vfxl92Kh8NCZuqqmsLmNDz464CXo8NBsfME/5Kn9OFt6PyM4hMeibwHCQ79ypLUTKSp+Xfbi
Hj+q2OVXWWPrddkZgqFwHhrZOxrLdiXi/c7QnjqdhTR0MMlZDcrFfloWarDXPJxCcPy6yEGd2ZC4
9xiA3tw5/ZfJR176HWbtTJTJOclQOVge/SkhpwZuW1Y841iWkmWP4JmgdI3ADoNmBM9IgXQPm2ij
E8LCqd37MpzBRPKp58L4sBJElOZe69JyHgzSJW6prxZAz82jyqJVLKb8wUFJIg+2bcCEAy392arp
7vVJgcVDwi0f4oyqQE8khUPi1TZ5R+S1kh4l3czw4L13RFaAbGKeIrUe+oKVfA39I12FTdG2OndN
902Yyb5/vYUGVYILoLTq5qFLIqorXq31RYlqIENPw/p3t2QcTG3v7dbHxLt62MEFMOLLSzhqOZYf
I7vWdhoNhcfdfYHhRjaGF90l2mCd423zlJltJQ4YSGbXaUgE91hlVHGb1Qh3a/t5ton/1QpIXBUy
UZ9EoQIQ/ZPIDA1kuALMWV7otvk/CJGrycaocO7QQ3KnFxVnZTmrW9HBaMXfEiwvrpO7zysYgn7l
muNXUuti3eXL+94wqfH/sqQ2gSggl0eWWyDAjlFXY2bpRG5/BcLuYYQhYQlz4Oi2aDe/ivNKVD3V
n4y1ncSPLYTcWhGpE23kusrzxMenjAXiB0hQ2m+4JSssHfuKiNHw1SoPX3aU35SG6rzszXKfWt9q
tMN0jN0xe2cAY9kweeTkHtb0UU1qSrHPLupeKq5kkPAKtc72HkJS+I2okCvMzk59aywSZ9qrmk1z
obisrpzDx2HAskj+mne2IVeSDYWeChzsWqzzl1w/WVXWz4RhgYvRj9dxfC9DkCKar09hgdMtqvRW
fAZMk0ILyiEkyVnufnzA5DvQF1h7/7jhoMkwXiCoE2EAEgbK46n8bwj3sh9ZY7fAxfcoOvkrAPJi
tB1O1ddKwkQlFaOPtmQw+G41FwzUwjMQBzMmbiAOgMbTUUtq4K+Og0nKZ11x+SuYe4FGnnLcu/cc
XM19Y2P0gUQRb0bOb83mX64Vqkzbn1oHUC9WCCenaFT57kXHnQFNFG+XsoN/DPWAcHJ1Wp0PKwxj
rvcLFzl2Wz0A/dfSeTM1M+Lr74wJX1BTkcdauHX6iwBkRpDf0yfj4h5NfMV57SP4w/0VAuCK0mGj
9o0qcETCiLS63idcuH8p30AbUW7/FIKBdNm99xjuJSgdeR5deYpHwZhk1WTEg+I8lgTYnvfOV7VA
Pes9t9HYmV3Z21Q+jsijYHbWdGeZg/fyHyjSOl/m8Mecw8tBJfwT1LQ/HNlGzB/CTHGX2T/QDgzd
GGCXBRMn5EA85ShZcJrKz4XLj+hjFk+gTs96hIEJuDrChiRZw/kvOC6aPcqkyDmZ6vo7MUatSZEk
A+EhsrdEh1FpKInaPIzjAgyrs0RRMhVzrawOAV9bqboGOhQ6YDGLvJOVpw1SV+phvETFGGlFo6DM
zZiZOHnsmFTZw+V4sOyQoL8ZUfs1Ynpu9geplIfTunYv84Mjnc8E+A4dRyqBaVAI8eujyRr2/EdP
4T2NZitkgMJtZnmJMRgwwVhGOmzfH19QnU7yHZas7Di5VWZ5BGH0UarOHbdnvqwekuM8W5WNUQS1
atxJsLFq8HsNtqp1hZfm4vQ5WZ+Yg8h69OeBYBfsfFfp0kICwhaeAXeWEmkK8qDjrhxaHTp8u9F5
9V1zvO4PvYaAXhzzWOCLEa6md4vtmyKq05KH8F+qwt3ug3rLPVF2QUc9R6z4/2j9PjYSkU55qEwt
MlRkR8MyZoUKp3I4d2KIopE1QtGWB2+W1gB9WabcVCtzSBe47Xe99C3duHOnIhG5m+3zCUqpDtaM
vzBNOpOvMJGnBnjgJX3UcYcSzzOYezojTtATPnGZHPnn5MuTlVElA2DWWCbgyme20Mm1WdXjORAB
2MPblVnPG+vyMUt/Njgbx3Furb+7ObnQPz9DEwpFBdjQnlx7nCmzH6N03KjnbGx4DobKm/Bf4iKg
WyFQ6+cEhXr6HLNWmoYlIT4wnyrLENWJg7bNf2qpz1/QilOtGycocHA9BOJIBSQIB2BfVlS0gaD2
13j7QPczWqtUgFFx0SIHny/DVKUhCxnhY6kwGlnPbvfYsEF/L5EcwFx+HR9lMUpZBWsIr5cbCnY0
PewA+wihUFKgf+psTk2mF/+HIcdhixn0Xf8Mn989eySCi/v8sKIG3fGh+TUG6VBNHYAD3Ej+JPpQ
7+mkHxM7QHUjCvfEUtTVk9N7JkM5kqTOZa5MZdTIx5xY7j97tEVwvJ+Xt2AhBrCE9Ufh7CyK7DmT
77/VK3aFIrseMB2CYQ12pnZSWJpV502TTzmllfr046uaRuGZm2p0/YUMy+/4zIMOdKJWtfHFkwkX
IVotf6YaQRhm10Alr/FvYK+dlo06t9w/5gQd5C5Wit/LthJJQ3UHWZSs3kcG5YWPsw4X64pPZ1F7
1BmCVrve/V6H4yKhR5hUy3ujKgM+dJ0uCVeansDpo/UDJK03sICm/idC3qoV7064KbOdCcY+XPpk
RMW0rP0WtKPbszJpBqyAly7PlSmAIrjgWrO5I4wI6FHCU1P+7FVR+xGI4o6tBrmRAaKICEJtwa9H
wbtLFVAPjqtV5Ag9CsH7A15T8ZXjI2EODCcgXbjb3FbLNCAlv0uIVUvrZK6fBL3QoI1ty8bPMTbE
G5i1zSJHnjwGzeL2d4vQBxcm5Fq/V/uh/Oyvmmg8Jw+fgsE6wrr2zD/ErtYNB4Tl4u+f0NBdvljN
+SnSl8SZNH7zrNcVhiNxg4Vty9Gg+ntHgY2KlsJFDkSnlIsI0M9v6ln4VIrWC4D8fKmuhLX5tILt
4KqQ15ePf38/HscasRwz30mEIxBWU9OCfSHiLyYYY6jqwhyHom/MZdOoa8jQnFfo7JCvhZLxTRKg
nZhgYSsiTtnY9dB/tqE5U5kvXuUKkNQKytwWOICyyU3C323at+eZPukgLixZ/hig8WigAnUiN3ka
/l/YRV4Xp2AvcGYYB1uoBsHI1HWg/5LuS4vOpbFyUvaX02eyIFZhssG45UyivQ4rbmp8eQNSm2oa
xEUS6p5FS+XK7ROq85MxmlVDfUzf/CHLtNOjU9nu5dGN0Ar+fRdagQaV/wpREIpLwFy6uXLDX4mx
VopWo0jSOWj/qPf2jvpKGPoTCCQt8Zya4Mp3CnqB+nTGfPVESa8XvNSr8a+qBdwJNBfIiOPfHAe6
zxg/CWH3q6SeveqBb1CS4X31RgBLSddcX7p1jsrRj4Vj3D+fbFC6+AiwM0tKLiFFcWz3rF60oOao
4aWB/HTJp03/dv3N46Cwn6M/hroEI2vcAzOxH39BBg0895mVHWyoz253gTNFIU9LQ8R+GHdknbmG
nijvdieg6k1cBS04wuXWW2+T/dfVnZTb/28cNj+T+3eVB8hF9gal7XzVxqbI6VvtnWiRhXDVkjnn
o5elVgu2D2s/uKm01cxNIF8/deu+e+1jYKSo/RC42Wm6dKM9XORegrL/ghi4Bfag6DM5ZhJnYbZ1
++3oVMQiiH43s/M1KgfQ1atSY4kYsg38Za+t7eHyHDUk2GHeXXTLo59UeyLqtBVqs1R2uZAEYzVm
kwWzwjXsmUk6XxCwTFQTWQZ0tT718kLIU2oceXDk7DFGznX1waSEaM03AEHE3rc1OlB3AIMGUg63
45PnvDYvildJZMXFLUJr1TkDg1TWgpP9QlXTuhGxwA1OaOoErYPNyV2+VZ4kS1BcPyan4L5gJpz8
uvjP3pTb9+0l09aDTuzeZJl49F2mT+uRW/s46DgQkPGWnUqNPi9EOntXcDPAxYikeppdj1vP0/Ji
+A5ynMW6OnEpNk3nDLsPH40D/Y8zGJRZXt+LWWJOHqMae0GkFUdU9Vx2HeZrbky+Bz6J5ncT2e6h
jwR7vifkcqFOr4PgbnFBOmKSX+Ug+mmbhlE05Pn6cMmHY1Pf6A2GoOV7JRUUJEQjvEolLtYe/hdB
glN7r95d7j+yeI1QN699wFOlTtUP894XZ/Z+nwBSuDAmODjMeAYDdI6gbPNGW2+Hu/YQrl4H/fdq
HNyJwkqGx0IL8a2XCnOweMjN6hEqZmmrpyUV3h7qDdpC7UxjI24CNlGRYMZ5o2c/EHFd8ifT4yf1
sVnzL2vgPRgamDnFhQbUZ3PBRRLTe2YH6QEyWxuE93vk/Pksp/sYqATvLguRVOU2ym21th9f/UN4
NZH4sOpB13RLGQbDmLmqoL8kVT5h7sAP10ICO7VYaAZb3kLalMgtcRDtFTxhSQqaChpdYboa9S+q
3Cs07nE2n8O+5ZGd84LINZCvWk6ZURS52X2UunBLYwvVEwtSWNy1vffOy1jxLj5DBjM2IRMsqCoj
gAJ+iU4JpkAMR8qN1Ltf2MEq3ocY3N+KrYU+0vOTnRQ8xK70ip2aj/2rb8lQt6eVdiKOMhi9El/b
ZfKGckZFjNoquGPlAuppe3bgc63lR/o4JRsHZwuP2RwXSJ4/+durS6JHV3LpnRlw5ump51m78HXD
Wnl4cilu6U8ifqQatcLa2CgomgBLNconRzbyIk7fukTSb3m1oNCzoIKteUF0qast6vpIOkGRM0ex
Mly4Mz9kiUAfa4Wh5yqGoBOJ8lIsS95gwfk2btjokC+Fh6QJw3j/Fkkqg/oVBmu+hSXifd17hdF9
CufmRNQ16VvaZ7f/R5G+5JSunDr2wHYzgf6wk9GP4Fw5FrlR0NhQGvwmOlXotc6kOxz43vMsbBqA
DbRvsM37Jw686iYj/qknFu2T4wqT4VXrfmTzdVHWoH3jtIKmJY1z/LOYUQ0CP3ZXOzw0g9q1PRyP
uYwJAAq1l8b0yjf6wr6lQTGZdYOZTsZeHbD0yomeEgmFO25XGgG+AXs5sO13LiOGyKfZFavKDn+J
zrn3/unrAJX82/79RmhfOaG/6GvCL5LEo90RoLnekarDUcSfMLy2sgjys8vrr5SkNs8WCTCihR1C
6L8P6Jp54JnUJI3t7Yefie+FVhZeX8f6VXfs1EuhwTzYGv4xB+uJhGc+owsWKCxi2COzAhSO+jNL
oyy9EfN2J8np53sAeXn0jsA0zutx2fGfR3zNZmQ2/c8HajLFTFd+Rm9k4jy4q1o16DWO/3/AHwX9
rTEGlMe+mmtRxcSrU2mGwtVED2Sa8TYpiAIS/t68h+GqP+pbr2W1fzOkm0jQ2P98rqd7Vblj2Gq9
wR80B2WeaL+NL1fd3oCajQBY5KgFkSBwCgRogjkRUA5uE1o/AW4WAmBlKkTz149W1OtlEqzmWBIY
/9vtuhgwYqugDGmzZoIpF+Ce5JGwYU1HAm+R1tceJkOZPq9VzTjjqFVFxub5daO5XX9zrguYXhzu
tRZ1EW0A8e8dzBsbVt4iVCoW/6MCaxl3ziRWF0UgLDLePDyFqzoyqZqKucyRskxR7x9ldAuyQB0m
+gqCAA4k61JzwKOQIvjcWGkJeA/DdwUK5XwBhbpLFEYGZuEKhEIlEuiGwXMT5jMsd02wqipw5/CA
jrYPg0vJjoBKi6BtPodnz1WIaD7UJZLYfcenz0u0mvJKxwZAQgfva4Wahtl85qlw/nswHVaWSnFc
dSNNnoOt9JI4bNo/03+wX2tDosTDZrAfNHiEmLJpvTTISiaW9He+8TAOLqrUBwBzDLfa/ROzFeDN
YdQYcftYxGiYh7p78km3xWBt0VdJh/v/sft3/gxtpbfAe85wvM8bzlGcovMWmMouab2B+wwyZrwg
D/GHcFD21mNXni6bOM0DY3a8nw8/aWb8R18Dg0UwKtUkTQdhG8561PsnXGFagoiVUXi6CWVEr65s
2JPqCoZG+jkg9HNcglYsOEne07tSiW5BReFpxB1Xuw3JjtITeSlmTgMVO6OgWVT0uMf9PXX+slG7
Jp9eJVVSZRGb9wvgGD1XGFzAcdu7JeGjoZ+VOoq1pmeXZYDbrewMh73Z18z3nm138cOmYNN8MJZ+
PFqQMWqQWdvOVogaB0tqjUMJGbBgsfxxEKm/h8qEP+PuiRv63VVjiv29rx9SUthzlWt8r47K4LCZ
kjPnAcCDugreM/fFqunOPV8uhLArN9ptNGB19+8cymSfdyIlb0lMCTOr+VMNU6m/pY+0CIgfvFm4
tFtqpGrgbeMJwvJJnZSl7tF2wkCEBDQuAFEcG1YGk7cq/gBTA6Wyp0HqtFgbzniduhxiCLJWLxpO
DgQIhu3aVx/cdRG2+U9PdoqbT2FW1G/Eq0sDVMF8vXUPO5WZBACZRWmDkjCywYTiFdHkQbU4LbmX
ndh17DqJj+THrgEC+8LQf3OLnJaGzWh162DLQrsxaQJ9XmcAvKvs6U/FQBAOqHeGyJS2DDr9Nx9x
fr3TIQlTAgUz131QiZgHbRFsRcarmiLLUEGyb+le2NEE1D93xMiiUfAbSqL2rUaSoVNus8VZzyzi
RitDxJv8E1ruH2BgGxVDeVUCtOb4zQu0fkCuT86lOt198/T7ULycO2UFSGr0s6gQQ83T3w8RPVt1
msL1zdJEOHEPE3RQIfNGuZm4uSakrjrnnvPX0JpMMBvrr/QZ1eLuKYAgcPaImbrTr4Z/6Sam6Jgf
r0hWugmE2iZU4R/xJQXbrhEwoAgx1+ylQ52qPZebhhwo1fXFJcnAT///7JLlkK9/J+WjCxU1rFRE
AKV2+x1cUjJef9+YoTT8N8ALuBKZDVyP3PqcnxaDGps0MqdeZ0zRvqnY6JWIonazEF8Fw8bSj5AS
PPdNigWfLqXAHJuL6LseAg4djzqtERGUCWjShtX6wfJcP0EhB9qtGQUKS4ueppF2nWIJplfOz789
9nXsKGjfM4LTI544UfZBItJDH7/e+z4dOqZshw7UE2RnBYyCfFlGVrUQ4eRhuqzZhfIa4TlK3X8h
JFaFeoB4Q/V/14N+C57ct+dHybiX83+7dBU+8vwhK6A5b7BffvpYSD7RpxKOco5vaLdGESI9UgUn
oRV2Swj7gDO94EBpw/RX8BB+uQV7Z7rM0g9bMxbz0lOF2xZdJq8bwRulSsMcepZMeBFUWcVt/ipZ
L5x3PvRSrP5L0dhSvjuq44IVtTmAYM3VjOBQ+WzE9Peaei/2rSw1ZTPAQDmzrMKMY27ru+d/Nk68
x08ZclELOrOOms8JJ5POyijWwZ22Tzi+quDETxMoajq906ig1+NHmK7Vajkm3iaOgQiiUk2f4nx2
GXPPd8id0s026jSzBpbG1SUY3Dr7nK6+sqMtokY83TLiXEsi/JmTcXaMj4jf4xM8Yw3XjW6LEkn8
h7H5Kot/KDlNIxdaG4yvBItiDpZ7uNA7i/HjumEYVXBlptcs83X9Tw8WXlpGI8jMPA67Ie3lN0Q/
0sfbJ+LU6VfnxH0NMPsVbN3GodNEDBBDsK3KTXTq4ncF+w+CuRu6OYxj18EOBXjWEhRZQTgZ6fdQ
dAi47M288YKM7XJDmMNaQ+EcbdjIOCIEJ115jlAKxLaUnFKWFDWsJCkc/bxQ9+oZp5NX8Q86J4JH
4ThQiNTGamt9wcz7bxZJNyEPcIi415Xwy4UHmQu27woymTFxQgx/GrUqPWSZCr1mOBRdiB9KBC+1
uLRuh8JdCHvBW+QLmMUniM3NY7Z+K8DshzzFR6m6XBT6lgoRVkHEUn8BDNnFIdpRH2VrpmKN/c9f
RxRyP7Oo0u/j8u/PuIQ6pdwGqPlvmZ10l/wvK2q02Ykuki0FL8SDW8ohIOBKAfNlKM27kdWP0Snn
n3c81QtKvb0RRzpcDJhpG6ItQ4U8xqU306aZ6Ln2gtB63hI6Vk4zrCKRKaqz5zZdIzBY7jyQWxEo
kR1IOTvHoMLbyi3petgQ3h6QNgaMGPvX/lseSl2Vk8a3Cml1seMb3Z/tSIvRThLARlpkpevwvQht
NA9/iJcK+W7hhXm2U0ahumSnrOOBbsBho7YxZz9LcZ3MquD8z5LIfNCBQ/FwX5SM56NvqrKKmRsY
1X9uoOdlaPx5J/fdrVCBHANNEY5jGxb1K9aBXTtqbNv8S0+m686P4weMwMWASe6w5NnK6Pj8uy34
VDzscMkllB+uxGtx/C4Gc8G6KF5C1+Rc0bx8at93p6TM1izt+yl9jZHqh+IOpUjj3BI8m/wE3Bn+
FN+AJJn5JAnPV8PVHKC1XJeDqz3OsdKeOJ9deqGGLstwJVjo/yIn0xmzs2piqBHUHvasQXWOM9hS
/pnAJCuhKfnbZxfAEDNxPw+R6xf1bP5h/13WaV4hi6+wOnEY/m1xP3/zNnZB2Df/PnlkGZNI6Qyf
WwWJhFmwOeXa/KC6/2kRvTweiv5hR37IDH1MC+Fb8FkSC6s8FnaEhmg6NCwDIzRGTzMCpLlT9npL
N8pcClp4Dp092FC154qSkwztQl3lQJjsT8jC4KzoWrgzhhYvzi9CPSWux4CmYCU2YsEfke4tlWhW
LJ6/2tYhkeUyDzJ+fdE3G6sVzydIa0JGqoIeCoKKMzmjtkPXNPHttZQ8ass/qZnmSarpg0ufs7X+
jUVQc7eEXDX2s7w2XvikJSVIDOIIRaPuWFCvIpqDd9KOi2nUcG5JAtfF974JI2xF5zGHBNLmVY6t
6mIiDteoKzqcPZcEpMq23MSGV5kh/VAohEhTRID3FBTmyiXB2x73UZJAHdRSHZkX1W3+PqcgBC/x
A0YpYRJpM6TSj3msJ9LIr34CKFg3AG4eE5j85xkA6D7VoOZGbDDz8/F/3FEr1csegP7Lkapivybr
5B1HfceAvJ+yrUATcmLXSvJsFEJ3zwWDUmTqBlKIQwzZAAX4YNo2rRo4UM/Z70qQc4saCi73W5iv
3Wi0giM3sp1qjJXI47FlFmh/8eDoZOdJEEYzluEn5BU8jDZkEW4EcfuuECXzrB1x3aFiL09LHpxk
4QISfFIvEA2L6vNRlcl8FwwkVAzl5rJ+KT+lijbl2gfJIEF3V4TSqObimpkI1d0AM4Ilh5giwUbV
1bXm2SKuzUq3hKxY1pU0zXJ60XZIZoAxcYEgeHnoPZ82dxNe12oC6nF3ZodCftIfZaCzqKY9uhsQ
xST2Q7AXbo/joTMzxBBlqiyyCzw5HdL6w8xr4EHZDVci+JCTnW/8TUfk5InpGUfdJNlkknJgUcg5
5GLreUpkaXCMkwhpTsMC5n2T6cRylJSPhGQZ1xJR7tiyloAXLlcyBRq6VxFd56FDg6UOJBI91oBs
o+53eqA2aOlOrRnyuhn+dQD2GFBtyrqd+Ug1KXkI1sKQfsg8n8zcVBtnLuyK/Fq5ymKMDfQ/hZl/
lP5e6vmFJYR4KGROYb9XQmherjNQGPuEVXVpT5GRqHNKw1hrRGXq8A72UzN/N+HkicPDrN9wiNsy
7N0lGfLVmST3/S9Y7y7aUL0FQJJF5b4bNa+exv4zkMEqAIRSuBlxXcScPPcgAN8rp0ayzmQDYDwB
P6+Knxo8afO2i4LhJ7HbIuZDv7Z3zyrA4kH6evfbkd5fhw1jl3d/XuBFQkLJzgHuIu2mAKeeDgVb
pmMBqFKb5paewJJXluNP5CHZAKpriUbuz34dRIM3899I1gmzDwWZP80+CFilcHoq4nT0QYwkqv0X
YRwATGLNMDh3htU6sFoii+nLP8LOtrZ9wtz6BUKHwtZrWPlnnOi5Ttlj87FdZzpSgkGiJYJ2LAVr
Dn+wFUwPQW7YW9ziqPHvHCCvRlScpjZgQN7lfG68pCJQjERPL3m3x8vYqSqfWLjOjPEZYQRlJTFx
1ksxHyEz80ayrPy0dg8rEZLm+XCmPpHQKAN8oF3qg9m0SFi7HkwUhjywKjMbSwlHsMFOgrYWYkly
2XAEOiythVYt4YWLsAtR6Ci65owXi2bXc8+6wI1JQvp3n6sql5FPD2rCZFcI2POmlnVDWXbcdNLd
OfDYlRY65B7T6ujEiTdvKzj4RFx6yvt7fwodpZTEDoKOKBo9euGTvqfBD08TnA+WtEcS3yeWnwPc
gqhG7MsR/YbfSA4eE3n9pWlo+HkzN9gZ51r/jCDW80NaAH760RMEQxDQ3/o7191ptsr9qo72jIoM
tZrTaY8+FzDSeI4tzQtXqn8Qdy/UZb1LLG7tU6bY0GMZyFXiioP59RHjoIP9+TkLUcyrxCzhsuY+
tyarT9juVnr8+Op52uXGi7Eb5Ui2LRq9LQ1jHCIn6zaKO4dRLYl6+CkxuCgV4rUjB13wjf5A/646
5IGo3ikeQRwrIy6KSO3XQolAAX1BfBTAqQDO7tTeuA8v3UFtRAsqXTI5BHab+UXo9RBJdKyVM6fA
JxYaguz+JI3NfQR5NGI/vVxmS/GRevsREyS9TbZ2EmuoizamBQ1xd6yrdGRpGNZKqSK51uwP3WJK
XAQ6as5FwEXguoiYt2wozukPSIZOIAGnX0LTW+NDyuyrtVIaoIdqH/sI0kWYvPpcuHGSnqaPtSG/
bfWuhMlxNuPk6i6ogcoZji1BA4yrQicwdSmCmZHXHfJU13xVE/pydpnxrayuNnjfgB6KrCuxKBqx
qmtobu3Io2T+2Dk5XwOLCdAZtY5e2Yft2khgs171MFRK8xIga8TaU8WdZfU94AFDDi65fTsQCzql
9Z4EIl4Eo/VCtUX7IHdybtHPIJvn9jDQOsFD3HfBOmQdW/T47E98xx/q95idVso1CaTBfZwIU045
YwN2pH6i2RwTeuQIRrjFCekjMfvzu4UaM+9bKRnXeymJlLqThWKX/edMsltx1OWze3Cw4PG1PniY
8H2HThdwwUjwNSuybHN2qJkFDoY9PGz2ZfzfWPxVJa3N0wgrxQ8i83yTmlRcfjwWs1nx1VOiLXWC
/TnLjb4JKczg/hjr85AQpfJ7uaN7q07GzID5T9P4u6ZFU4I6lBQzwxYzbEAj9dV1GqG+7bk+T3G+
B1k293cmE1GhafgEf+v+gGL2GWFH6G3dYB7XaBeyStyrI4mRYW9t4Tj8JikrRb5zZIwiiydmVq5a
jk9YNkacvapYzymVsRBqTthcCMpRE6Gn7P0omz/VbGKHbt8Yc5VoxPFY7OjeMu8jt5mLz2UzBJOq
lWtSrurUOZ20m+mjIBmHgDJX2jT23XbhvEvNi0ebcGpbxoPbLYro78ijeMtDsZlYUrdNsLxuDI5u
+3ds/nB3Qj903jkU8gbLhic9vsbLVOlVj7klCGXb7NLrC9E08Ely1LfWzyOd89YLLtUji1Ly6Ove
4OVy7gcnyOczMUyE1YLj9vr7DRTSlHo6kkL3fWbvO253DWC3RhHNc2fFiRTyK+CtCilg7HdKI31D
aCgaFiS8tI9pL6u9DSEq27fdTQPvpbF6S3sLU/ibvP+nW1FwWqUnfdvxXKMOJfWthSBpMn8NkgFP
h6uFvFUMwcfoRkYUzt2VZddSFhN1SKmq1YEOWyDZWgFNu3hNhdp+PdXsPCv+jrQWg4UYfSlMkMj3
p4qom+99N0LMJTs5dSP99mw0ke8BKoWcHN0rkm+VeqgivKFhF0e9bU4vibkpjOB/putkolYY9gU1
poFzkSRnr8j2l5huVSSqsha75qiLdeg2i+t8YsFFjkxO8JvCCIhsURD0mZVb4M0RRKSU98vXJowt
3N7Nvc5AtqttsJIgdOP5+dhhVhRMu+g+rysmSqRcglP/3gTH9l4BvqMuGni60D7Lky5db7AfK0Dq
wR7Xx84X4MhK2MhTgAytieZTilsz9YHBX1tdWxUIgL4+NhopXuAXmjedE8t06zf5/wuXGvGuKOsn
qwzIAo3+w9NmnzWxjqCVC2ypOWJPe4Igk+dq8WjtTGXlyDZ4mFvBZkFLLhkzTK01Zj0QG+3Ap66x
ndLlIQ3O/0PKoSy+70wMrUl8p0q5UavAis0q9OxE/oVGcaznikohQLc51fiwDDtCnjmt54OMUWSa
ZvWTeLbZ3oj3dpIGjajE0WUjHyV1ZmqTb6G/HZzOSduROdm9ztaWfXelze6x9r1P1nAtqv+SoErS
4aH01ZyQjgF9rbe7rq6s8RgAcSyfsUiTkqFfwVYHYn+hI6sp0GLKL5QeJF+NnzbZBnm/RfAaRQ6d
nxB4qv3YdDs9XpmH/mlp+56PAu+srmjGmib32Mo63NoaZRLNhLJU/UrcevatrlppiedLEdfgKDfI
M42R1bo1xq8vJTyeubftmI7sceaDsikc3qv15pSgyfwinMZDj7bKkk2TR02ALbmbICnDpIT5rXzc
DRVSHAxZGxUl5uKE61AqwEnqd0UAH1IR2SKaTwCfr3sBsPN5unxeISrViPlp2eNsgFLxubSowHK5
2CjPzYYT8kBNCYGTTyt1209hfE+4lGBe/YHF4hM+jnIlD2W9NKjO0m0J/0BkYH/xXX56/3N8tJZe
kquemf28yfoKppPEVCcdVxjWhUBGISGGae4WEg3rhT8boKsSqdkNU8TDmzMEMyyFM8P70u8NPaym
AHConz8ZWr0BtaAZDmh7JpgsddRsvSYJLQlJeVCZ+afd4fgWOWfkrrvpLhQrwv1BUzKp/fI3HzJ5
0IHeVmlmbPx8lDgpQ5ZF+rUA+z0pw7PMDdbM+fgZ/zGK3k7wbhRHEm1KuB4eX3oCJT4Bh78LO7Pu
UqMb1r4oq77g2R6SIev14QBG682nU+PffJzO1nzHlKPIOYF27Oq3XxFVySups9R4oDUCCATPLpGl
Ot/QD5dtZ/q93XoIahaoGU1WeYMFOiFGf8/xfp8r0xdxHq9QmO0dKj+wCuVh/kXNWZ9G0vxzgUDm
mhjywGiFN86itQzopKEpPikJb0ptVMDmReqO39SfdVs4kNOGr02xKLVEmohGmwuv9sETOzMBhlX/
lOTBrI5dZT5BmY4naj3ekNyZupxUF1oCVjvC02nAnSCrc6j6fc1jvEemZjog35beZKjeouNmzhgu
kYnD4ULm3+SwbbHJ7kfp+KIhGl8w92KDfRa+6CXXlAKZooDJ74aKoBaHxBny94Uad563BzphjfnZ
+Uj1K0I2NE7w8b3TxhmhwMdaDtPy7zqpqUhyK9mqJ5gYR5ws7JmyUhZIb/y49qZft9yykUwHDYvd
FQUZ8pOr3cgRDZMEbSFCOR4EivaIgt2s8h9ucdNhYYzOS+Fhr/AlxlzRZhmZ75gPJ2SZ062fxCLS
qmnVohuBlkKENgIWhkW0JPDqCcWVi2hS4jgoIuZNqNLxW58l3Xfqj8ErUHZsDe2ZuBplTDZuvoCz
JkCIn3tzLn+HxrtyqaxlMzBXV3Si6D7cxj3Va67x9JuJnYzpXCVDLL6403mPzK8qLOcpGBb4zJfS
vblfkkFMO8t8MdTl/Z2CAzPqWu0tURBuuQPrrJYNVHh6Xy4eKCuId7V7DThpNiuIzo5DGMZ+sVSx
LtkIG6skdmUtuyPR2JoiWR9XeYFQwwhTgSdgx/2M9PodBmxmFtoB00MYzUdCE9LvxmYjG5hTzDIw
pUHsnmPCrifQ5iNeQUaBm4VzZFqIlSi/8HyXrQaxbzl/3zgcHj8WeRNkyXERQFB5GtgcLmidooDu
sPE6UsJA44HA0eMsY41Froi4YTF7kDQ5hXl4KGTz7r0RONvQMJgn2D8KDBz3ep8A8TKcE/3alDaT
2Fi2RuLGxAny4vZVhVMUkisU8aGWqtVAMNUDzhnHTHsvTUfwjBmkQjWiQeOBzCP2HfVY2h+42ELe
MdvuGQGRZRgLUmQHix02FnNOWgDUBXYhHU4kMxUmFrq5jyHAEDXiVbXUre0FGdnrNVsgP2gYraDJ
jaRbnUDmUoY1i8p1nqXefTfVtuHSWRTNjFiTLuwMIx4T8QY0r9lFjzWalT/rAMc/JlYZfeY7xCHJ
/EskqNJk0E/rJLvkIx4wMmcHKcFFnsIjJZNjToB4Ig6VpKhXu/5AqgaMrPgvmCjHlITwzTJ8imbp
vNUK6JvoEpMEzPwEdYWGWN70cBMib/z0YZf2i0KjanEchKKcvEiQ1aAnyiV1GdyuF4vgsP6CPTiY
L7oqCMv/vT8xRIGdBa2chFR5TtMARvCGbjIDxjd3KkCzuGynjkk2HKly1FvrpU+O4OI7xQVE9ggJ
p1j+onbb5mYlg0NGm/zIxmp7xnRmwFENDCkDy3kht4nwJvdHHBJ66o2g2B5+KMkXRtMfwcUo3oh+
jw5EHz8mwD18sOLtPCuIWWm43CVekhkKFE2Ni0w6EO5w+rxwuoxEjgA2oAYIvLGWZ0VW83TQ+g9z
FnYnPMO6SbHmUWqA9aZLXSobhuuVu1vjNgybCndwqErkNHnvyRQHYJNvpv9w7tJKD1/YaGpRtMLp
qbpmzu0QnVytrcJP5FNKc5NKZzXvSt/+3WXCsMtlUKUwxGZ/7VqdH32Jo8d7zHFKr2GrrUL9kqY/
HUWcc6tH0IV+z8HCwv9v8bqcEKc1yxl62sM5OwLZY+Dals7LPgaR0gqvL9TJxLRBroMt18HGcVA6
TV29/5qiqivF6gEHUZJmvsNcVUuxFHD8pGd6UCToCJ24P5Drh9AjbVSmSAag8Av+FMWYb9hBx2WB
wHYg1OWvTDZcxYcaKdBY47+gdAZIcAHIs0Oiqu+gKHbFtACbXYGH6iz5Q6TuJDbITHuSGsENbFHG
aEurtxY9cODp7/B7/4UFokDu8IDI3cImz92mgHcw3ciR6+oXi9n/7q/SOZowF1HpvkmqSNuVZ3N/
zhqqzM9Z0hJtrbRVJ9mPYh/wUqM+Q3hsw2y0DbueVij0pWSAUHscwSDY+2SNtnaBBXr3zFz5Im/Z
fGfAr1x88X8zVUeD9Fhx+zxyQP0LRK64C6MYScl7vmw3NHrkH2Q2XapEBsKEod57APVzpMpTKJf4
Qx6fQ7Pw3HM84v/W7QFXMlVK3makx3M715+sKcHN2GWXG7IWvhLvc96amieptjg2M6YV3l/VHpDm
9uydikrUJcu1OUmzshn4jMq0tNo9rywKBaKz8f4dbNIjyHibIDOO5DRdEQE/QlJelmSqf+xVmRwq
NzueqGyKbgpWHPou4GMddBAmCQkCiqYb+ubYHz0oRhqLG3aUnSixmCPzG4V9n2Azb8yAIe4xDC5L
2o78KvgSQIBW0N5p19RtHf9qRcKvoCKgXT997hzN/6AN21pwS/GBjdrhjX/zUN2O3iWqnzmo3TBC
PiOoMDde9JNPfZJtYOOTg0Tymx9TkTI/EK08ID5bx6ycS2cEq2zbVGI3zAjJQchrYscQpBI/X9VY
Jyg6EMLGhyJ0BPK51QPpJ5Ea+CcezWy827PDLdj/aXlLNhk73HYKC7RrhMgUMZxqlvxx3QuGXZbe
DWERu7g0o4x4x4Q/i+UVwdIpzWlwHcvJRpg6/yjzepRVRAhQhLA55wKnMHDXv6KvpUVntSYq3fS7
BQhI9Pyu4DlCtDZjX1YkltXxCGrbJPMM1boSu/paoDtu/EciRHX46C4UvRYImJOwy/dMaoZ8y838
McGZQd26/61zlzow1vZgiLcTmly2B2n/6ToiuOJ/rdxvv2dt3okpW3OwcGddlaMW48I4RQx/A0l9
oo1zgnj+4LyPezWNyqj+aINsnGAetFlE0w4OqNMrExqrlsGTdU1RdGBu9D737LjMRijAge78fBMt
R395yAYYtGCwoKWPX/Aerdv+cV3LHbV8aUNA1BrpKKhzSedQDC2uR3sNL+9wH27JOe6xqEMIAIYn
m1QGf4eyiapXiE2PkUPEikH/SRpKtuU3G/SEUqrIJC/gWwN5O79D+/X71lj5ah7U3saAWzPVYmsF
eSzvePmakkF61+A9TBFVdByrTbrBP1iHtYtWD1S963DSRlayq9U5MhjPPpgYhkBTLKBT22cntI9A
1iI+W3plZHPrFoMpiAkjpi9tuGQQmW0La7f8gJ2f/zoyxiXKeNBynSKLTBInChzKcnFSUMgF0fMy
ifDPGad8MqwQhPJwG1ZuIpACdX1+stkQUXzme+MArdx6xTTEPejPIEGx+wdudjL+LRe/nKXiaijh
WTPzwE00ey4HDjYqstxfhMvFV9/C5cjnQ9vEEAFL4tw9D5hihNjcm2U4+30n84Kl2RZaT+4o/rhA
/610zbtS0VKJ2IGGImMGBJhqRVuBv8Ani2FpwCUmqHtX3zEPg9qk7dc/bb1VzdX4hyM9EAkiIDL9
cBlzUhKhG0fmo2qDTpKzMxPkDY3XA4I9bE8enRrEtcLWhCqMdrjltpgvMt5tA9Lmd3AK7+spaLhQ
QE/3c0fB+lWPfXYLgtE467bvjDrBH7AicqCMgitC7qkacRnNUR523bpygew95575bjP3rPGHFoeU
O9UScJkUHHi7iKa+TvLAD4b+6xnlVN4OGEoRQFXvba0L4OFTkWpHDGW6g0su0sO9dM+7ew3LQVUV
RLaLt2vtVqLtyd0XIzmn0HVxgDdmb4W42gxFCwQuHXfRWij2HbFFzRfScx0zipB5Dpatk0FXqp0N
ZNqGe1+QZeS/+JOenk3Gn8ZG/6KuLrV/qN0R/FTmxy7MFtXy8lidnBja3AIoEvWmevb9bkHpKfKb
8f0HRKRdfsrKxNauDX9L/qGhXu1AmCfnUPcRvR8xgBbz+lgcwdFZ+Fhu1SfNmYVVw7ttBic+FYUY
MU2IzoXGQk57yhlhtoASWG9Sz5zEu3mFiU1mabVQsdNBGDkwcChlDR9KNy7vqLKFWZoKwYBLN+am
dUaGvk1PG8G9E/PnHn/ZfBjVYi6Q0mf9AxT9eFmwjqRbIQFTOnGk3gRyXoIucy/kocJpmL+OUa1K
BDJxvBg6+6xUiasKZ1Ji1rdTsB8yihjoQgVFm2KTWhWtoBwxvm2HPFu5ZHvljS5zAk8z2kfiYRAS
U1Yjj6RerOUlB1cYr06Br1nleK4eFmkasg6h/QHn3TVzLAf5twOX1g02QrLmHe+eTiP1XPgSC1IA
OpFn8vzMxQ+IaoF13GvvVQiWHm2t9QEdPnd0HSa/NX+Afo05K4Hv0QxhidhMmMmkuYv6OzYe9akM
hTQNs1EMbb7hGk8xJ2mxggq7G2gvA5kNd38jRQeqNd/ZICJzCvmMQNuNog4A7Ps4gWAdIZR67uxq
iYEc6glV3D8o8GWaVdR4Uq0ztOQYGpbp8pVYU8+w8fYH63gOkj8xAwYVzIHpNCeAPmxIPjgXtZle
yWA5poeh4+HZTB4y75F4kLa8G+i8xctX2ybCUmSIuPV38b8mnqg5AUod+aq+Csh86rwPQsjDXXvX
IEmemEwOTipAWDMRHAvx1YnFMEMHJ/hPamOfZ60ydthklzPpxrGjO5DG7KGtCBq7fxk9d+kF23Mt
vePGS7zZwlKVbISSpUW16D7lolihhZbB3QgOTQIWEE5/zxSpZzOLGb3luW3ZnvoW3dZdubK+CddI
OYogvwkybmZVeIH7YP80ZEi7dqQUawUW1du6djKXctOZMswXJZwoIwlFCqkLSZIk7N1O9QzSrfkA
SrKpry2g+y3NFiW9EMKynLSgI/G28WNhsfnO57NLLG7nJmOLFd38hlxLQM3nFQTfuH3pwO29jCOy
+OtArCgAx3a9/RD5abF2kqNcuUSwJSS0dyDyZOvAtPPgzHYraGMouf6eQAAq1dVal7Yh1StDv99b
ShqQSUOdPE5hw0BHiehGbaoz6v1TDAeZPItwmrqwlaoK9TFWxy6ftTAGkH8EFQx9CayBkOUisags
AYFg52EbOCMg4JvWn3qjC/LTF+WmtZod7vo1VjSYk0gsroeh46ycswYpav3aIZJvdewHoAmMoReu
hcM6ByVzKYPR0EjUH7aUHO3NeGu3xD2949u+IBSZFIBZHdOIGs2SM2nw/78lqUqeuEnGeTA5gzRs
7d9aj0XsIDSyQUlmX/5yFevf6yxcT2UdpE0uXiXXhP/cyEw589G1dJ36TCfqXcJeRsRxTLgAwHdt
rlctraNOlhMxh5Al/EG9THkw42nqVZLB0OZHiuMllqlEV4sMfQgawkU9sgw2bOzD7m2sVpCGomdM
hGqKF9exX8fx8qS7UwRvnoltjW4eUEQlHcUYL9WG6Sv7lFNh+NkevFFGIgLdJjdjnc7jl2dMDDL0
3T0spMJyEUFQKtpD4+Oa/N25s1+us5/G6iNYqgkMpcrQIZF8kTEa8LqtCraQgpqVo3/RQ2McApoR
MdGoqvxIueviEEASZVPElTWLaZGlPKlpjU43y4NdZEae2btAytptDkzRy+yFz3goJGC1wcXGI7iC
jhUfUVwC9/qhY/1/l1kBt8RLJ1Tnff6ssxFOrm6Q5PHQq7wS0cMJXRb+9x59KnU0oSrbzcjb2Vi8
4XxXbvxisvL32/LksxVtIQ/6DqaQ1o+tlZZ9H+a2kFf+zuMabmB79Kfa/p4YeJr6bOVkLR8nNXsO
z5irMIpIrCA9PyKKzafFkn4KbFw6BcmxUbKW82um5mh6wL2ejBcd6AXaGxfsQ/0qzNYE8hi7mnj8
I2nLLFOxRFqZMUh/qn2ikBxmY4E3EVmlQN2TaVRccMZduu4o5pQkrP8GcghOXMXAWJEQegzinRhm
b9VdqVsuLl8jw4zM3FiA68mp5L8mjqUvUM5QOeVOR5dAPr01OShdnlWR9OFDrOfJ5RFyHHiTZVrP
I1C2nxPzYjdYsoTtRbo4aiGnrOsxiFYTSslnGI7a07aMVQ/7jCPoWJZgwopm77cyL+3zfGrdtgZS
ts5JaE6neYC9tjZBwojuECNDLxFgUriiohFbnMsd4hrCrpeWVtIrKkObnOzp3y9StRMn2H8Lxosu
lrhzOxpvLRbryihWHZLeuCPqKiaykzzMJD32mOK8PyOdYALWubjzdBIqC2uqyUcFyQrl1Dk+nMaY
iqjFwqf9vc7+fmFmC7qppzpwQWmAq1EEv1VND5eh9iQ6jwh38ozC83zid0RKc5c3XBgJ7xfpCeOM
dsRoxEENWDnC+1AG+L7TBTPq9nvTmHEJPFXnhQnnRZ0cMO3TMoWIIHNoDqeM3LzbT7gUffc9M4/O
aS3z0WXMIdxDgcCduRQAT6Ggno9P69+4cloX96fzU80kJnZ0HmVtwhAhyI8StK/jDHskU7lwynhb
lTsBApq3NdSy+KgwZVptupIcSqdrg3K3zpssFa9nPxsOmunVaRUNysBxbM22u6R8+MMpccVHr/E/
58Lyi8f626Y6/p72KzG90KS23pO53bq+jq5up7IKJoly6IvC3Y+kKqHkesUx5ziYWWr0+dvbs5Qm
3X+XFXCIpksS4gIeA2y1G6oqJndN4/4xqRiIH8moSmqV8+N1+spaG1W3VfOpS/eLtDbmrj9QW27Q
rF7UcCxGdIcwuSwyGyQqm2mg9uzU+9swY84VRiugCKTdi8jdHs4hVq7kAYWwTbgFbNXvPUjRDQEo
6dsmi4TqP8wPgQhHMwLtIWkmhi1o6GYYHVplbVGQZyojJWyQVr1RkL7zuVqJ88PoCmEfcpS1Ghp6
oIt69yYDrxdrNBlGXzjMD/HfcAyyD4sGx1ugqq0HXdDufsta9uSsf9sUbN5y8Avbi6wi+Apxari/
RPvSQZ1aATtEjpeLVzDDF4oesDFr4Cj/ZXg0z3Ys26Mp7KMeD+R9FUpq9Z33p3dkFvn4iPAhITOC
MZ87GchPlNVmwohaJTRYKDokUgJEWrBDWVbIL/SdkXgBzOAhy04nWA92C/xXfc05KU+ojuPbnnAi
dqeBgtcVKaatEgKrmGLJWGw7sWAkoQBey0LqHpKjiVPnovdN71OSX+XgPNW5uUjAh5tOFr/8Lfi0
yxLuteu8aThQQB8D6ZC+wslbQsT46MC4feVPEHynN7mgJWQcxg89zKDr5kFXYlz0GtkYsRONkucJ
suVftekGvqE/cA6vSrL7Mj+ge02g7rh7a7Kf+VzPgZDY3ta4CwDPalY2IZluIvK6FIA9EcOuk5Dt
AXFLnP/kt0IHyC35Os3G8To5Tmy0egr+StVqPOwSrLPCrONunGb/ud0qYKf6QeJ3R3n9zILaqZyj
SWfOAa1PYgx9sOEe8lyh7DVVNUEMBloUfdIk2O8v7BaTzGyfAe5vT7zjoFdgXhB9g+5j71Cp+ANK
tcJ7wqj/G+FZmt94N0S865AXw5xpqETExwjlYc9/nK+r7R3IAxeHlmFXsefvzDe1BE3FQnrZrF7Y
r4B6enZA7x6oySwPgbpZ9DrHOToCr7NMrdAlvLY+UHfaqjPZnWfgzjPO2Y5WzyobF3CkGL07NOju
wmCM3ZRGJo52Xw3HFI/A3IJRihiY8OpClSOimBk/AWREWpQ9vVk5htQPVOENZi06EaBJrVGdxYhc
RgaC8fd5cuDwytuveXgzs1MBnZt0OuXDQnE6IxBSiIFlmtX8JLrf00VZ8s21N2ei8Blv51fSw28j
u29di4yvzy7WbFDbhb0sXPSYmXCEmatA/IVn2mx/7+hdn7HQlUJ1soIP+g/FdV01/Ysv79frcIY7
8aZpkKbAx5QiTxFWcGlGjBEcEYYsjJN5G2Xtw9qhFbqGEvzN47OkgjHziI1xfUAa1/z7J6WBHuR3
4yY/4nRBaoKqDAWjSkvP3ZUXU7JubrRxIiWlWMIs/9bA77HLtqJR3HEoEA24ru5afR58uFlHhnje
GjVssmMo2Mc+N/lZOHhUYlYib2lxsMQhddrnjheWgJckue8dMZB7seZs1pkTS2z4E9GxtMfiQPCC
bwTV8OTfRcgf9QqVhY6nmicAriS3YVUplDYoKJiDHqdcYF1IzpEfwEsQZrKmbISqJ6oNxaCOHDyE
RlZnGogXDR7MQ7fRcQfPE2CAhoqVcil4VSIhTjDPu0SvwgLRwiaDgAw0dKQDDbcxvMBMnEaxmhA4
YA67Cv8PsfTn04F9GIEG7Is6HipPRbIH7bXiNGhSha7zYANTQ+qVw7xj1MwyDDI9DRHGWgFWkXqy
bpnl2GX374aaJcDR8GGCM0ssq540nttifA9H+KvwAtEfEaYkXC6UmCCsFEiHjZutyDwOj8I5jrES
SfJ+Q9FNyRy4H1V94OxGC14rOPB/x/KT/jKkeh/U+XP9HBfzE8R/mR6MgqfOOa4NXXgGU0mjsW3V
BSESFvh7NxJsutgngErm3HyM5YfMJhrWqSe3o0QOFmXTHF4StHFAfNAGwcKLY6LNQ3ONULsiEHIE
givclECw49IAkU/MuYgIjHxYA7lb2PZs5owEnPawG1lFeg50edm8cIq6y28eLY2mcIBrI/u/UR1F
WWwnANn3Z1btjfSaGv0TAUwEiW7FQQkeYWDHLUuoBU8jbwmEPwRQwMBNOyzTo53lIsmumAwFz1uH
u+q+8AASATzxG128avomLIQqPsaVw9ujvvTw5d8DisHQWbzkfm3jEorBrS95GKNALEhhrW3lCVuZ
hDAalsLMwQc64hmJQgYfw9CTonvimVl8TSy9lvTFyC58XRkznom3QuDEDya8H5r9nzwl+CSTp0Kr
VtbUlOYTKxIPnIg7/QlLYX/95bo7dMkPh5iMXwhGpWEYusmS9TsJbpiTvtiBfukQhtrwNVQVKz+i
EHPO15YR3kBQvUTvuxLwFV72VdHNKa0LSfxLxPFHA3hE1fSQZIAHe6Sh6GDpAwz7TfANvmkWsqWO
QyTlaVgkjmtjp54hi6xgXnGRFhoqy6Q+4wZKE3BDaWO5NSDj6pQrAW52C8tLebK3ntOF5N95teyR
vG2mApcX1T3w5J+Mwv2Czt2ksjcl3qyjK6v9YYwZYgN8frgyZbbEgWbKu3qHnTDdA69hWcJykpil
cqF6HZ97RztgZ3GnHGLrE8PYCGj1PAMxpl73XUqtYGL5bbewFkip6+7VuoZWN8i72aPhpnSthWgJ
Vj6SBXvd0ZruDK4epGd10QhgWwy4z8xyd8vZRpsdfHfvaH+GTNLpjS8cgxCm1mR7OGQePDuIGTT2
1/qWBALXpUZ0xCoPFp5fCgDtyBjFcN396OWawsvloONyZTmFBMWIQ/iC4GvfVC6tbwnHMtP1z7/O
kHi78C/aagthDH7gE0zcCaYM30F98fYGiNWWBju2ew15RhXhhtVSqxgr9Fn4J8o/tgysAOzRjfya
PrRIRMgJvcgi65Szr5UZPW6HlVbka1/MrMKRdMvadHVuJap3UbLcaHySVv0lXQhpgFCFuHig8kvp
WvFt97ci/5QcevF8PkKTyQYBTfhVJprasPi5rqrMtoaFp/DYjaF5KS4D7UqUpsEcpdmdodlT344M
kojQdsHNNAeHZP+xOv5jSOscwOxCYIsu8FP43/GGE7gityWL1D4vPVb0ARMtq8ueUqKNDaWmulLE
egSwQGoGHX8YhhaxZ2LbGX0Rvs4TSoO4R66+ky1kncCDQMjKqPHvyzY/UnoumLymKlmX1wh4Cuii
kh3dYQLYB8UBsGoyHPF8L2hg7XG5LamlunbgEUxZy1pZi+h7RpHHu1T2e7B5yepAuE2bviGe3K9J
WmGRf3A5LdnGkoZCUmDGGj7qwockNWM3ZZ3sMNt/eF4GYpkiZHrGtb1sjgvnp6HDRIZtbb3wEihm
tPOuFBKfhYG1XjJ1VgUQ/lKJP4r6y3iqfkc39fo6vZ+Z4bZr+GJ81DlJcl7+qgs4Z7CKXMk6Ag1Q
QBLoDP0ge63MAtDHYw3GCNOrlCbjol2XHHN3IzY58zA0ihYlMCwFcwaRHWzkFPFBkuuH0mhA5T0l
oamnqwvKpK1AyFoswndhHvPVUp+scMvVlhExFKx+GUqMDnI39BUPK8wHdxomy+rShiYQ2hgs+GQo
MB8RU61PUlcu+Fwd0dapnRxF0+IY0RHM5i6XRQwjAYoU6PtYzm8nsHwrhKCoVkDWAiV8uGHiorQs
BMpWv7STbdto6nhjJTMBVXuc/eAnfsEUlOEwSAzDGVdzrRjbUwPmqMCAA4WtCsu2U5h7O9r5ZLjm
1/OIGSL7DM/t9JKKXFlU+Gz6glQTF1sbCevkBvtLSSXPMac3Pxi+NYYnaQRoguGRtUpPPFYo+bdY
2isZ3PS+JAodr/lZx6Jwbb/DZ6PAUJKckpMJHoXVrk2e8Deg6StngOjvfqoKkXDoRSK8UlcPIyPa
IDVT3JlAU/jhF2rzXK84unorxed0xZdBeAJeBSXbNTbitbGcoC7us0IEXrcx8uDxE/o79T62CTIs
xTdNLoXEbUvijYp8b22pGLx/pfu+/sul3MB1/dNuynPJ3TMRqsql+IjAb8+qqU4zvH3gyLJcnTno
C/7cMS1pyUuHFGXnI3xU+PgsX3Z9Y1qgVtOMqvRauLBSyCXErDcb6C8T9c89AfyCa9Os9UvHpxsU
AFFJB/dy4T4uY7SCv3emWpPC8hN/I88kp9B0dsmj9Uk6mDU490K+UdqTpbL0DsusLT4d7Lmr4XHo
mRcXTgFl622OE9ytxCuWA0actoBWY51S+TdXSjvE4kWnm16evL9q/R8GFOqxzZuTPvEXc7i9nHXi
1NyWIbIP/rZklZUSJHtjQh7Pg64ugnbojozs24IFVWW29U4cg4FfW7dnyC+NhcyhVdCi0bfk1ViT
cSC2Ycv9qHNciFMoIZPH3r8tM8RNrrdmLIOFRtSfVG+JQmdOG7/SQeZDCSy3WnZdv8gcAnG5yRfD
6gnoP8nfzWtCcOoT9nGsWdKrCnQjcWSRJjJ4cO35hJBx65lsPvIMWTJifkTTmBX/YUUVxjNYqzVB
y3Idnv8cOiz5AqkqgneFAeEsZj/u1FrImcMAkeGUEnw5k8XhgdY/iWPEnf99Ynz+itlKqH8Wskop
SQQAxQbMt38DIvopmG4D0tokA8hzZ9iHWaDgGJLybh41ZV+JaBNCPhMExEfguR5G8Wo6zlPTzSzM
igX9BJ0VZoTiFAGadnoNo8gDIqLQiNLoQO45tNzxJSt+spkOTVMaxo3NNmH/GyibfFkvlMgMc1V+
zzrKcpysP15tXpMLWYtnwXZc0X7/Hz+zP1EPI3e536L67qte56109j6DyFes4llyOwkWheMfn6MQ
LFYrf+maaIVzWcIRytOmpZDDgaPI+JBcJUuT8O1p900yDbWF97b3ZRzsR7Loz4wNjod8euBb522G
E8ZtVh/I2dFO6gxMMNizd+R9qWuWc3ML0rBC2d3U71+o40zlAzZpcTr0I9gm56DW0pu0ld5wTCw1
vW8451n1CIy3dm5lyIjJbiP8/1JBgEWZDSAhuXncH2MnwdXU58h6/tRRLW1vVPJaxMBIYTScBMyv
naxgn7jChMo1wUofsw34P7T4pLh6E6CX/efnNK0sUaO6ALSAFdOZSqrfx93cOlXcSGDRwmnfafmE
Z4Kx3sWLhlhSAMJKd4VLDUe7pCPSn305oFKzcmW/wOdiqcFRiGfZObpZTe5Ke8+0Odai6hhwUHb9
VgiEr1hm521xSxqm17dRI/EwQxFy40zxZQrxhsm74s6CFxUIhS8CGAWVchmzHRagRKG+PL9eDnEb
J/MVHJnJ7m0pVrZVICGtlzSrUq3vDPuvq9F5aZdn2rKWVjEX/MXNAPVIdJKMYmp4hStfKVKCKfB9
0h5cOytG+lOlmVhi+yQJe0sBD/jHFhoOXApbBqiOId6ooF6uA2Hm4d66eFC2Dp6gVIMS+mpvOJJL
BniGPZ6MxNCw1Xgp1FNmINqFOcBuBpLVKViPYrVDDTjY1pPgJ7S5xlKXeVV/B/2MNKBghaWvq0Fs
yburqOVPY/eRp463+3vxvxcMZLNQgk8ktxNHecG6YrLDvL94r/oceoffKvnd18m1t3tSNYqNPcRs
20JTtK6UynuOhz1drWugp/FFxu+wp9cwxUPMY3iOXtq78AQ5HJuqsxLsxX9kYuqn4wVzQWMly4wk
7Mjkz1c0LyeZbS8/zXfG0ZI2k2hfPjZwXatkeKeqahPzhlgkWUa46AeMthdQg2oMYi0ElrvRRSuH
leq13srXGLE5UzVFxK+QwqUxoCe1fXGvl/av0UikkugYyocejP1Thr0SDRYWuqZv9LM3HSKR4/kq
g5mesN/t3c/H91CUBfsBan4bEO4UNnhS+g8Dq+AUKA/Cux6D/BiAkisWHalnUv/7oi5MFa7h6z9J
wFju+Gvhr4BFnmxTJ41hbcPQbAsUGwPX2FIXzKBeQ93vLjchjceJfzRE29j9sq5pFNwSdke772Ce
J1eWuJGumvXpaCK5OqilBAKL5zKo1CTaRaqwPZvObmxWxBhUeCSY/40feEtNSy0smpum3ttcrtwW
b5zW4MZt+eK6RxgqquL4GZLdrs4pndX57PyKhdzzAcaedei+iUasXm+8dWToXr16Hgo/4QIeZp/j
bGmxpkrsJI+BizKMuhjnBBn3Zj61BBBvX0+L7Sw4LzFTUFs1HRV6XtT5qjEzWFj4cPo48erpMEmg
XTUvSvj6PuKNMP5dJP0H4CCQYuwM6jGRuUJ2xEJoNxfeQ+mvO2GQjtAjOJ3uqhTCPouSuHKKHA8S
htnkzWulGF+5QRI6uxbb8GSTussVX/2l4WJBVlt8umEGFmHRAR9SVOpOHDc3DveabAlxCyMevvkN
QA2kHhTICy5QKgJk7NIvqQNERQpW4hJdFKU3JBP1h9BIHSQgMe5ijHinq15x/zlBPAYJRXttpe40
S32ON+zsc+VmyouOSYtkuxcjXL+/6lpXY6NIMYN1rKJ1cfD1HmobbYhRLykRNI3jsz5Uvy/ounjC
pDaKh1LGM0449sLUySva2EZvafFxh27lKmBv2wxNds2GPwbrU75FqAz60knsEh1Fsd2ClWX4xjRD
0ikWzhPiXKw4OcMfRZED43iDgbDug7kWy4JmVJuwe1XogsWHEvlcDdmRtSvQzEHDiPpA2Y5lIr0G
OIppj6M0qKXJvk0y9GtdpHqZTxUxS/2V9O20LzK70HA5dpPXu39WfVVNtK9l+zavx/KxBvSiShA7
WUjQLIkixl9X3r9kPPKur1bgtbbaGlflzyfu0vc4fGem6cc2QZJtkNny7tp1PJmaDZS6S9GlFGtM
L5IOzSW3ulJDo/LyeegfSDtn39mC+7if+/vYAkUI017EQA2DPzIrZPYst9KTszwoexUDrv+3oRcL
9fVklTqjPEa3E8e8RSGJ7iyMdaJ62F+C8h5PfsE1lnSz3qp2+DYyK106sg0LxZtD01n11eiECZVw
BFVdpU+GdTiyvXGTR8QOxGNfRsqO0joruhutpxQ2/knRDyxh1mO8i+Gfl0ri7Bpn5SghylnaEIyM
gwC0G8iwvFBJqgtNiA+YoMamX52hmmZEH2WaR8QNnam2oFIXaaLsRpr9mPzlWkJAznp+Ow99b2OY
uGhNkEFUaGQkZN2+TKLDhSMZNcrP2uFd+88K2wM2F8AcbP6snDo2s58Cn8/YlfCmvNhF+2Ctm6CL
jCelHxsvTxxxDQsykHbOzKRyiMzVIo7r3zzzxCVQf6B/eL6MpgYcQGCCtIA1cw3nYlNL7LE9Gtpa
s1vN88KtbKuKHqgi6sQJDLyDC83w6M27jlLRsrT5eV1RYBTVzzWgDRpRiG1HfrweYYCmqzVf2sFC
fIKbmjs61p1jcuCaAFX6YjMD9x3df+a+XvADGgG6kDIaCRvSgWm4/delyF+7AZf55OAmB7UvCi+Q
ma3j8QyIDmjS1mKDu5HlvtducIieSJdqg9+71jVSlmOVO7OY40qvhzP0whuXcZN5AfE7amjYL0iD
OKtqA4DK17HBo/Oc/3s/ORuYBXp3iHaBEVjOZ7iACuYrM/QkhEvSA9NOPTWO8QCnRR0xBDALD25B
bkpUyGvm09DghWIwWMFEw/+TVxUrlmomXSJxyKIscDxElsP4bZVJY8+obt3V4+p/RQhIHnEY5+g8
X9bm2SASye6HDIWc2MQ6NmYeso3jGJPSnx8wmrq7IYp42ZvhgKwjzB3nVMnexlIZV5Bjp0HwPWsV
2OoTM7Lz/9+u3DLTMcjrFzCPSsMTke4YOXFbOArWa4HdOwlFDmDpK/HYVAd1cY7QevPTYnflo6mW
wMr8zna7Q/DAr9qKaBVLWio7vtkbk68YxXWkAgKnC5ueMegCEPAwlRdLFo9LT3BBbGSKemXbg+RZ
IU2sJCZdDpUFcYqXWix0SZ9EeqSkMhq5644DQliq79PNTM70G6gIgmq2Ra+5zehPXv/pNr9W8IoE
tgltB2iGeA44JaU0SCk7OostMV4Fv1gG9telqjOYHtSu2ooOCsfGXZuTlxw2s3Ad2JfDzSdjYAvD
exTGWP3PJhAdL7KdbaHOaLuo62ctCucJty7tfVAXrBCelFhUwBZoQ6H2z1MDIPOdwUq9xmXmMKhh
LcctuSAcqWavAITf4PQI10S9b7SLk4lP2j+oCuj4m7z1uTlpSIOG/R0QZmtwROH/uDCywTJLmqOa
LNtMeP6TmBmQsPU2JSkAwDj66G2ZJfQbTjcCY4Ihi2TT4jW3vqJdc6/EDSnq96w+y1VXOXWiTRUs
kcQ6WCBQcgmR1ail3ub/yK7SDhxVodOj5mMHjm7nVj/AJ1VbDhxFGCOSfSV9aJ+hW9b7K93AbGwC
JJ+HGAa02Rh7v0KHMmEo6wAgu/MKchqY5wPAcQhvKeC7JsMn0PpQebc1CRnikgZdVMGwhVW218Mh
Y9vB3FpIwXVMQwzSg09K5DJCLlDESQ9djZGR0Es8JhH2ic/Pr/aQ2jUHY/faqrptLCFhKHRWPMss
6j9bDFSmvzmm+qi4RJk53MYqNIyUwTIm+w7p7Xiruq5yRvVVJJ7wYF/A5MpJixLGcvSm85tDO4Vr
hp8+lHW3ROuCGVsqgRrXwJVXgNHUaCDnbj4phSehrElD2UW1eT+9HH2qyVnZtUU9Pkx24ePX48Nk
yDioUg9kHR75XrEghVElGxemWrnoezwk3o7XG4KwiSXq+AUiifBIi8xq/ewjYUcvYs380xBx/sJL
/Jz3m6+pYDGEJjqA1IrrogP/HNDNjtB/MySoI8N+UMXkJ402qm4uVzBYLi8fQzSeRykMBgI24dHq
Jm3mgllhVR6Sdss5BHvf7kdPx1m7Y3Kw39UaLpmHMLc0jENfXKmosRGu5vbULYJpCE52GKIF2RDI
dX/vEhqvFPe22JwKA+2CzWl1199qvCv4u6m8JNLdRQmCG8FiZLV6hLvhrTEshvYsURtLGe8lrzBJ
CfPMiKLn884qPNh81ncutNTS0BbYS1H4Fp6R4GyY5nITfwpvXr253duCEVrJRbieKM3mWj5YteGt
DC3iqwP/2OCNkqqi0Y8qcHRx1ynh6ECBvkGKLiQX2kEfq3l0rm9UDoJJ1O01KBlbh61dC0SQ+oS2
bXWIE9v4AiO18H+LRGUGmN53o2ZB3OynOhdlUrkV1St+1oWVoxE99D5ykROTaxK5YAnABSpyQ3GV
wEUYhWlgcLs4vJI//OdqjWr4igfdsBNOHB3Mm0dhzj0sYrhpdROohGD6A0FRmg6B5wLfDr58blxv
nc0IIVTbfIu8ftuPBqTlakRie/1qj0zok9FWjoS9jmzBnYjspW+MSqI8IaqFlsthBHhm9lRxHFZB
XnE7vGVuhNUrQLg7Va+QgCQb47CcMt4awBi2dR5T62LuI5qSKdzBUK/IAxna+1iFMJ9HW/H+2OFz
x4XxYgyPTbdTRTD4OtWXhP9St+0iLU0Vla0thWdpAGMqlUCdHELULKpz6lQs4MJ4Hth3On4OevKF
LA9Tt9sYJQtG0PfjY5eSd8sp3dCPgihF42H6w8UCVHxRFUZb0pRO21TXNHA8i740kBvfZmnL9Bm2
WBYL/V5/AxA8Y8B1nu4xlgzbwIZn9OMVqUygIs8N4RAs0DTecvkW1B1S9naL+TUU2ANZmHsS0qUV
kIlg4j30oKb5g+UbY1u+G/rTYnEMJsal8LPNA1YPq0IpA7WStwVW8L4hD8629CSij1nWBvp24LyF
Gh4DVJCFWNuUa1WvjUVo7CsXwtFoLVA+l1V6AlnBKzi0dk4pXaBjf3VdzCTTs5eUlzbLD9Kn3hqr
3Vh+w8qYBHjOGp0XIFQh8JJXpV8XxHo87Y8JslQE++ZfgHS68Dg0j1JaKjElUorRk/wUmcWySOFt
T3ZjzJTAI/KcDEP6A+snDiSXMYv1k/X92ciF41xuG2jfMMR070+hK482YG92WLK4KhXczHP7hB6F
XtVrt8YjrvN8MVqGB6rJvHnEAKKr74ojakIk1DmNefheTqm2ToaqdRbmiXQH1kP2ThSU4QZMpElT
00kEYURX9SGOUg8m2dQeWuR18SzOvQSsOpugbWw4YBE3MdcU4qDBz6e9eBoBFEhY8XnfnBxBVAdQ
6gwyxC8Rfic5YdG46HYhtGj0gMd3jInpD5rtsAqXtmuxaQUgI164OXLv0RDDnqF7r7tLhnhMjOIR
W/wdgi98KEn+oUMTfYcXjO3YAIfBlhZmO8qHQfy63R0Gwj55cVSbPd8g4o7aDBYSJ763T5ASj48l
F2nXt6F766gPgKuoBN58Y2F9fywmaYyaPwpOruNXd9Af/RSGGHPSzMWCvVb+pYvysZI0R8cn5lSn
Ony0Rch3VZ0mQuPDyA86ddRg4pDABvWI+POJVJXXCJR3xxTgNf1HT+Dqc5t5jDmhB8qTofGad35N
7dM155eVFY4hEU+L4rmP462309OCVdWhhgzmZRO8OA8bxLbTKL3BhZfhYPDzso8VIF+Yec15feQD
qzlLEY2OgMGFRDeQxoh+QHBwpUg2WErUFGe+6KvwdRvrvU+YioMqwg8kEgcsa4hsuhSK5jk3GbNb
8j/IVpEYVtaL3W78nOwz18rYo9L7PMvIQtKAeLybQDw5cB4XVdmpZ/PngqOegoBmapMjVL4aUBD5
Rq9ZDqr9h+egY7IkpQclWFIq2gGaItydtcFK0U0sdJ60oVi7XCE2P6ykAVw9eFxMIMQteeUD2Hb2
jqAYgznzTIHR1PUWhxtEf8FMtyzQMD1xP9vyLF8GXM1EAm294EaxCKaEU4yRJGoXin378vJL8vv8
bHcc+G99YmL0aDL81DwD8A54sIS2W7XQpv/3LWxbbJIgSooVC/AIpr3NXOfnyeoftIA8810hX0VU
Vj3gqzwGa34arsBVmfgXAkE8ls6MMN2plXsnXTNPqW/2qz9G1pC1N3jg54mqVcKD9tX74bFIdoPB
AWSFEHXRnGwJZkSFwaS/EuvctZakgA30b/9yoY4FQGoA9M9pebOG/yuX5MjJ+bLzQ4FiEMJsTCiU
V/LAbau/UJEmp9YRvx+2kxS9Aeum3q/6A5Y/2lWdcyNfXaBnfMy+CUSv59pW2ssklhF1VeXk/7j2
TfxYiNokuDil60Y8NNaAIzMFgtawfEALyYb5l7zqZwmxReyXpoTWZqSsx/mstK1s6+4W7CN3IlO5
e3nu5h/N9/Nbx28Kq18yDBNQjlZcMwRgcKRd8+IR8lXr0cjyW2CHKgzNPVTvguRB4z0syVRvXN+I
DfQ1wP7yJQxh8Kaw08qPva1eoOXhy6Eb2OZaJy8XFTLpErtQ+WYmPp6IuXPXZ4RONSl6OcXGzRAn
/5of1qwv2ZYqgCCCMEtkc/rUNkrL+Kc1SNmHCUau1DIEHrPNd3hxDXrPLr1GsiDy6v+gmBxRBpTw
q56PVJ4DtBxVsB4naaQNCsftERCnS2ZgQm3kgDSVaNJRBiGVbaywVFbVpR0CHA3z3tldDgqg2mB7
NQgi72KhIoXNZg4PGw5EDavNvIavqiZo5YFD+jgxctrsYC6eagYG/5g4RVSuDvnENYlS+x5tBkbx
NtlXA8nXft4EmJmIJELMnu7lduIJph2o+YhS1X5ZTIzFYEg9Q/57zqCL0egmO7n6Q7bdthadnFGQ
F9u44zRVbLVU3MiJRVHfcaikMRuuHfZMFOW+M7piwyZ3dDN8AGSbiwzXiGbRhnQB4G5CToVcm7WY
1hoNEQFstZZcLQZbttYMGbXtZu3OiFRB3pSB6l51wb/qgrv3GKnr3E2FIdlwlqg67GW2llyhLzUY
dEqm3ZP+hj2L7IbEqFEyqZ9b6hJhV+zdm5D26c+cYWRTct3QzeCy/xqYk/pYZnBU9mjmevoRLoxJ
MEj0dONqirUKtkjuWX7B3tEDBnwPLzEBEeVUyjmhgyh7CWpLbwXWrqgdUNisAYvmRsIbE8sXDJFT
dgk+qbWI8hxLO2Giexi7ALQvDB7VPXAoEv+D5IDO+OWWe9p8O317jQSzpSYDJ6QvVVxtZOQ3jovP
sLrW5OUNKcgxXULvxFN+uuoC1fCXuw5bIIQ4YgQ0B8mwhAtCiVjXQVL+O8yI1X7nL/JueoN0bXsH
1SKYuS2OPjIimJlSM424iKU3FaP2FcoL1JvF3r2SlnwSLjF0P3DmwJRhYjaOwV12M+VoanZxA+O+
pzZpJ4DcaY4g3EtKEiw/k8avIbaPzVg4KEKQlxc5AQ44y+3FAHfWbizFi3G2RgVwa0ewGc9lnNVu
s6JehiX3oOSeSqhfmcHevh85dEi+09OMSvMHscY8eafNgb11DZKUN0CCLKjVl4yYj0szHpOz4h/U
OExa6xPk2ywyJAGsPu/AEE+hI/4TzLdcGy1RwEySq/IRaaH8M2D8J2BJ6KKM81UlDrT4JQWVztf0
TdfMm4zv+ayVuKL3gsXJvdzpWaf4480eiOUSYVYMRzJucbd4ebHYaUxoBKnQ6VZYU4DU784ZqKsR
6J4AQMQ6Rg5ZJ4XKn1/nfIZ+qSoHuIhvPXRx7SN7FSnLg1Xy+Tj48Fp2UYQ44Rwx+XXrzLhwsaYT
fhSD1GhxSr9C6IDWs4uUI5+S7TrU6ciFV+mklPWT3Xo0oRpixu1Np/fCRZl+n0iglzxjrfbBK1s7
1nAT27yRJaXd5v+jEcUqDuLKIbE3gvnOD9q3ZrcpSLvEdGslIl52z8r8IveEWt00a2k9GcbfrJQv
3K/x2Ikf4pEuLkgDwDqIrXBQjuymAcRsKCnM57Y3yo5RbIsQ/MtahFHh8MPJfqAhjRM+WBcSHvQ0
onhLCBLG3w0XjPZA9NvTgGyE44QLWmIkb65DLpCLXE9TBPOIMWsZr8Gh0rNF0IkUtVj2GEPJCcOX
ci0ZtozREeiEXg6Sg++e8BVdYPs3Ig07Ld8LsDu4gF8c1oRayFCquDkhyJoozza14QKpB456ozlr
CtMi1UQwn8l5LuySOpZUUNyk2DspFeQ2PJK2IECMb0TThIlhYekKWDkRVg19cRg9+7n73DdVftTi
IVtgJduW32+5DrvQye3VnPzMvE5KfDSihSaIm4IlqEAyma3lAibYehCn6V4O8wv2p/IJEbCX8pMU
iNttKJ/yiGGSvPyQsgZmD9WFpNvy7JgcJ6NwDifff5Qj7aCYz1xEL7RuAeZHJAQkL7Gh1XfthxJa
QPaIctSbdhxTsn4OvTmp1LpdZzw0YuRMHoCjSh+j6JIZsSyoTndmfNuqL/O0cDTrcjyXo7NjgjpX
V482Tmd3ieimkBRhVCdRTMR3G7PstDTO0E1ddOblhoPFmUu4eRdTJZ2i/uu+QALLQMxyMKmje6ki
hxQC70FV6Bh5BcUn0OAxPsx5lecYMLmBCdJldgxYFbIYQ6RIVDcFUUlRj/qQNmn6gLryLawwxHZa
Ehor8cuk2377GGrHNy0/Fg+rNAvNMtk/ti+RFO+ydsPfTdxqhqIBoXPfeR9XAFKN487jwEQ6zbVB
SC6CYpIj/xT0P0umhtVQ2fNkzEeTnkjXJfT5Rt1m3WUALNFZoG6A+5AKZa92y4HOuY2Hg9GHiRB7
a2oZPKQdKIicpaEKHzeKkA8m9bB4v5PkA0v8OjkD3fRDrtIkr5N+osPPaDH+ZcI9J9bI1S2lI0PV
yFZ9AASVYxIR7my2pHkSeGI/jTg6MxWNuu/Np/RZHyvrKBQJflBa+2t7Pz08fg5OtYuG1+KVNAsz
xlTdOsZTnU6gcxsBEK5zlm5UlHTzAwNNoIT3MYNwNF4na5XOJ8YY1nYdL7jmQcM8q/M6zXbddRTZ
Ztnzmtr/zxOZlV+3VoyxBsWW6pfkQss9myKfOf2LbBciKa10FnJwJuQGrj6wfHbKKWssJ0ET+gkg
H2GAY0ftTYvxSr6cyoPRystww4i6FWCqHtlHAdMKtP6JffFJibNLX5Psive6cAvEsohQ186SkEEi
5Ljp8K9nJq3XDrk73sejpilFKMs0T43iInFVttsty3mAH/OqaT+/75l1ReL8XcpfvWtij8MZXwCR
6iCjo1Q1UQvuA2wNNzvBTP4nj5T3snjXN+qioHtlwwjG/9+OoEC9XJbML3QiSd6qOwEc4Nu3gSYC
WopFuViMKbYl1yG9OmIjirTuo0W5OLs+5bwrIlsY2TvFWMWsxNtbFjnZNKtGjdGy31FimqFCRzp2
KEQIzXrpyPMfIwbn5Hwp0HOdPHdKen5BmdyT4mPpI/a0EY2TyXAgzIJFzB3BzT9+v9bIpdOgbpBw
xUeXBbfR/sJnERSCuxm5z8sWxdl6wAkI3QOTutueN9MHBp9uj3di+UZo+PbeIVHKF/Ss9vEb9ynw
QErQB647PEHMqI2hoS3UiQ9MjiC/8xnqF72/mQsXFm+tTZ70recEqlaFihzLFwAF7BmKssliDoZh
+robvL8RkW46VX3NjSPgxWYR7LZ53M26NFpfkrNlZ8P47X6ri22uFpgxeZdR1XJ6edTEkUytsPiJ
1aRj+SPfYEwWaNbOfeihP5fjY9kqbszDb+Q5IyCE9bNMP3U5GuVnUTAfWKQiEkJicjXtt/CraK6t
pRjFOvCk+oTIdgmkrM9QMUA9gWc01acY1pCpghUFr10brz2SvzE/rHE+h1BdnqR9KG9esgFaCu5/
DeBsXGGePLYSzH5SClqE7nhKk64R9gWJSGG2AZL+RNdwy4m0BtZbKGl0zyl500DG3mptLyivNs/S
WcCmNS2DuLklmIiHtZ5Zbbk91M+RU58L7s4tzlYH1t606QZVpd3dZAfqT0mWSzkFnobR9o1kpkIp
JE+BUaWfaee8jRivjO3D45MMKzk5I3xFZDJ2CHly3mUct4x9/dhMNK9GkxREKmBC5j4NDdCplM+l
9ycFEsrL5Twfa0X8iwYcHeCKZVOX81hTeYl8faIFyGpe3hbcDbRb/2VSdn2ricD0y0PFoKrwxHKP
BTkFBDXjk2sVc5mUrRM8fnEu9KKy+jv6/nzHfPRHPccFjSKm86SUhyDhEMwqlg9Ky6munO070ZBh
TXneA1RrbTqg4gaP0Vxc3L3wPNp/Dicrrk3PFi/ujgiXyAwlCVdp+94gmi6QSXZYpZUEf5Ut4x54
Po8br0lIUXN0V2BT5bRQZ+AjmNaDmWmhncF3VteW4YYJkp52u1gPSGWpQt0AoOwM6w9uQb5rHCo6
Idi0kikaWXgxnAEcCM0kjgQ6Y2KGQZIyw4nv5Ta9cTQMrFV42gwOs/iSXtRPyxIWRpbbox3+irli
SmxVPQGJJrDomN8XE4b1qtemjHyzLx833694zy7WBjCNF7oQ7WDgtBTGY5w0VEe6aVaSGPSvG3Ft
x62Y/1YLkDzXR2M6aINHvgAikRh6q3KNqBysH4xTBgnK/9V4hpCslI3L3N1cAU0pJqXijEr2/qWa
NU3L3LXgrJT0XQGAAqYKUfCbzQAfsBk90XlLy+zEmhSp1kjHGmUy6JQl0XkOW0hnCiWzP8piq3Y7
d6TYNiNwx9XBip7svV6gS0G138Vj66RFmGCTmvSKfO7V4n/w0zJs79pAWyLJFJSGWvtoYDP42Mk8
JRUMZiK6qpy5FlqjzU8t4ro1ZhfQW+IxdfH364WyYxNPLy+hr1lN/jirUKcepk8nvZlguPJ/zHui
MT9/JkmaciHQ3NwQ46e0MfgfEi5pLjwcUsN1uy6OkSq9ET8aPlCOH6dtxuFw+Kf5gGNrRXOBQUWa
OsQWDp92H19JOAKX1JoS8U6dXsd39KHMYKc08pGYjxfSM18dbEkwscv9IufXWlHQ26D0w0TETRqW
HYu6n0pfuKxN9wmd6Qws5pJ4ErKfqX9lsV/qW9ZmROhNkf4rBnBPF58UyNbLWJQtFAK0wS+ax6Dm
+kqJYMquTSMQoT1LW0waf5nGWbLOEbghPE9laixowxSIgNT+jrVg8xij1WPET2G4bPFqEa9QZDoM
t+Qce7USHSAPihUDwHLoK4kiI5w2N+d/9zpFltEcRhGJgnxFXocxi1WmaBcHRcjLqi/NaJRz0BA2
d0XjkLebJg45rpAyxoi9xpVhXXWWIYXV2CKU5Im4MO1Wm1fY+GO74EGzXQr3DRQWecuA+yHALSff
yY7+ykvfG3pfGWTQRyZtLsqf102xFmuUA4w3ZmG/UhuMLziyyMfQwiHGo6T1ZhcUj7GpA/uPgg3x
BhKtg+kKSMPbtm81F6uCf6HXM9g88lEZ8Rj1CYikHfaAcJxuK3RLiUQkp+3W38BJE2xSTLL0rD7z
rI+/GjYZidJmRGW+siYwg8Pi4JvkKitKsS6VI+jWqs7IlC/FnHj8CG5ADyjze4a3hyNT8bBE4GXg
C5wF81MH7OnvI8oYZ31/JlzM+t/12ELAuW1oa8FG9BbDM6Mrvml+ivhJ6DRl/IDZX15D4jMNuuwp
ESPD8uMEYqjz8c8tAt3Mex1AoIfBaub+2WI/gvNEyvLFBJC0N581GlNsYWZl8nnJm3zeJ/yCGiRx
kKuz0G6/TAmRcb4RbHYdclvZlkyeGK105RXAxqXEN9h2cQC/9YMvDYYXOqBM97VEYOqX9rhb+Qdo
LUyXhcrLe/4JTPAF2pXpdZb1j4lCM2IcYmR7P7QASLhfyg5lyAlnVDpkzUfyuBVcmH4HF1j620pQ
Qo1qt45+HGZ7CfMWfiQ9eUQNLxQsgSdWhEbgm9ubG3WhDYirlvyrZCo03gzvp7WnEaSOJh58RokF
yp0OKryKjM143dRAcIWrn1r8C74DKCnhO1JI9YigSJ2pMkY3zWg9pRBwkQ+T7yzcEV4MxUGpY0Dg
enDyZV9/zpRzRI9inyqk0j5VsZqGRrXS39ga1KcgAcAYtm6nfRDsWkYC03fPk70cN3C/ufcGoY7q
MFHBQUhVHJee5e75graYCRTm1Wr5H3tiG0YfvkwLIt4xcvJuBlndllJSt6NVX4QywF4uywtrorUX
G71g7p8hSVILJs17IilshG+wNzAs0XcSX+jwteiC5pbpWZ3QdchsJ8kNnFr1Ys0rJmz4I4V9oNHo
fKbZH827af6NGC4uT0XKa1c+4bDuKNKFWvZCyWxboL58cX0bjo6B4MNqz+Tgd4dbH7LO2mENnTcx
WMGuzDx5+694u0erI2bOORpPbxBYe5eliK/LfUNpbH6J01N1lmevv2XjrPEG5/BTbrPnGqv1LopS
aZyM7uW2qfrrau79jk1hNKWjHzqj00IzOZZIfn6X9Xu/VnXsKZiv69ltLjY/sYAgr08EJLlKwDqi
SZBsxJn97EgXt60Y1eigji8Y4fR0A/LddTtMwoR3V0zLReF5FfhW8Sj2bhPHpoAqSQdSHemV47oj
nzF60xLnrtuQVbi8o4gf5+50nWK4hwZbz44SushzTi8zQkmpN/ZiRQt9Wraki7/Jz/vTkCCoyd5O
FXz7hFC15s+L02qIvPkMBYBmeYTl2fgHoyCpUoLgcnwz5F6e1xEUhkUOsJGaooF0jg/D2SMIZllb
8aUNOSDtf6wBSrg2PYPi2p18TjGl17lr8sHO1BnTvFSlHww0bOkYz1eXhvD3xRXC9C9zPw5bYvHc
RdYZDQQAdTCuZ5yJJEGl6SpG/lMPWRD5MZmO/XUqfZ8/aCOz+XYBNTT99xILRcM/YoehuVCFJktw
Mt3HxcifMC7Yue5pppwBWlnxvDpls90TTbafyFLP3LoYcdyqOA5pLPWjWxmC+krbPsQxcRVgPrid
eLTx1buk11uMVjwDplXm6SJgIHyxZ8CvnXmCORwe18PX0uYhUZVQZSsrQcOPwZz387XkjkoURVi0
y8K7S/9lwgUL4WFM7RX+Y8nt8LbHMGpa+Y+AGnJY2Si+S8lTvyVyR8YzgVLMeYdCNNUNJpEJ7NAU
5P9vEBulnpSEe1m4vuQAZyP+EfCuS7Virx8l74rF+EujMkRqbFs4vdQlzeIMfD/vDgrYEdBv7S+C
fa+NRY4//XSVkPOsO5JiqQHQrBcBnFnRoTH14Tw1ccClAzb3jRz5vIYpNw/b14GMsOhKgMbidAEN
yRh+x70FKK2F6dcYh0vAe5fKQK+vDnO6wGHPaeB3NfM24sB3yaSOi8wvGAbTmFwgY2xrO7mmFd6/
3YPFK5VYE1OWM4QZddetfP7Y7evPNv1mO+rea20ZTz1r+yG8am/PPM9D7Vwy1rWe+rUHs4dGJ12L
u5fBePsoc72bSTb0WsFAA84T9Vq3ZAQFH2XFZnI6EisHHJ8iwjQtXn04JPh8vvECFk8Ls7/8ddww
lkcLcQyqMBQTRRTzrjdiflZy8QDwnuAh2W8RT7QeBgpGmaN9e12WAJOzDCUmniq6GBz/tdd+RbKw
okxZyi110pk6lS43YXZvjmA94I1KkpQOB9eSw15AvZpLzupcRrpZBB/fANx54Rb6mm5xdumCYpXL
g8iEOcLvqfBubpNgi/vV0mAD1FKOZ+sF3kt0+KjVUgMVDPsK85svg+RJa14Fy5sjUgIABJ/fE4TI
vVLExaYQwAwsDrGiMb8HXIakrAdj7Fo6FbR8T2A6NykDZH5vhnFuqv+/KDuili1BRsfMe2Audb3d
vUcGLvLhN6fCRZ5qBR8YHzm0xEKpK8mHL8ZJ0Kv+JICX3/JQbNvXkAi3iicp2MJ6WJqFNXfAsYSd
eLZqR8SjTF1UWXloi52NILN3IhKczG+j/c6xsIFiVJ/jy1O+/ASN6EonAZwftHsI1QR98SC4UOKe
htzKhU5BDHlSK+99hdSIjW6mUi/sMVT7fP8yJ7gpeQMrrmGrDFQAo+y4oiKNNWAxX8zQ+Zk78j/8
xC4Zf6Rt5f7DSbY+BTl2XwSZkRSnKiD+/Gcb4nFBwWz5dEF7c1Ej421aJpSeyvsNe+z1Vwdw9guF
JaCt/Q0zPZnTsdZyuOoBIPGIiZelxl9Tw9bO8QR9jMdTg5a/ZNVgMYUjjGbJillGBige4cuccWkj
Pp9F0v4oEyIHIoDs6Rax+5iRCWMxKfhXCizkODaDLq99e6dw35sE71sKW1Ftb6sv1H1YuBwEFIwp
NVkohoFxNksrHhGBfRWJSGQSiXihXvxAbc93f5kJPzzzG+CFjXdG+U3h0ly2ihnOjRVnbMK/N/Fx
oTJ6KMMJcrtvrjErZ47ShoNNAjc7cwFyZSJhKHa07NUgzT24bG2utjWx65nl/u4562nuEadYVuf+
Z3DCA0mMSFj2rt5jZZWMZxChrsfBkJPWg4Wl942PTjqgpouWEDXpTGoR8QktwRNLZMkHpKhLqjBF
V1BUJxHdkiRfd44zqeLoSBc4umIIhHQ1y5TxkmelPbRCZiSfBUgQn/6lLk+6EpA7EjOIJnevMqey
7ER0crR3AEfwQcz1ed5Pi58U57C6R+MfXODm5DQ/feEARZ9ZZsPl9YwMoO09u4RL6gy4CU4pj4Wr
ja6O+liujy7gO1jMFQiHpCAXgDcUFFBWgjTcujMk25UeTZRRMVz7cdE7PXNj06JTQ0oCNb/SwkZw
tVpEFSIitIivEBctr2D8vlE0MxcofxNXbie425IzyB5MfEPTOxnVTDMmDPq9GgtHtpWBs+6Hgp8C
vgsqeBuWuxeodRjt1ojcivrODfSOwW67Y0PE4Ec10LZ/IJaPdtwpRYGoJkACapFmJMIXox4KBZE6
Nww2pDIgu86ZOkpLHhAa/rVUvNnjjku4Lem3ex1/vxZAamzmaRLLOASMEaUnEaRpPPBWf4wQszvr
asLBGyh5HVbKduAT0CU/E7tFCQ8Eb+5uxvLgCRi+90rgWbBDqMqpW44JziCoOiGFQUJ+nKaQkN8u
iKoHI7Wqbb6eRX35gCr7YzeYYaXUaaiA866oDzIigq9Ih/DmF5ONhrc/0AphxGUidEuvuuSrJi0i
KGF9mQY+EWJsuzSwWDHL3M2IbMRwXBsc6uPIQdQUURwfPou/1eMUxg18UQqWizjsElQYs0Wih8S4
xCMxYDQI3wb81st9ggskY3ElEYoiKV6R6C6rAaErPXImxlF8in5MB45+TtFywxqwNIOyI0g6HwYW
lEdDPvg++GvjAO7HxGWjOXt7TfbKEf5IE0/b1ng9QNtHj8c7lUpCAShGh7i31oVXMJy37ksYbqJh
fJkRTvLNtVW0LzkBgfvgnNWpJmQU1iLLWyqzIEtfyc9Peutz2MRtkVHiai22d33n+higrhBsKuZk
T5nRjoYseuvDRv6qiDy2cgkW9pMacGbAL6HF40QO7vgrig98cXMbQZMqDFN2EbTakvcwSUILe7q/
3ATP/sNSHFlSFFqStD6g63gXxsblyNH513ABMhvU9wFcxlm2BknqrGdeobfiIsf1l4YxZZ/LBph8
2NEfeR4icHueL1O/VXKLZeLuFGXJC3ZvkpYyEIlBIV1EwEAhldIFM1Ag4Wdz6pxUIEUwhGGCqMNC
5H7PdMWiCjGDfY7Fmb+MguxBhSq9bBt3bwC1hoqzlu+P2LSqduFZwOjnF3fGIXG8NRbXQye7kUtU
x0cSrt/4DrA/ppf6w3VmPD8f1lBUoCiJvNPa5+InKkZ5juSV0+db7QGAoP3VUE34dRz5uMl+I5Ai
z1Qfg6A6iTmq4pOIc8jRuLi1+hAoBjQOUmFjD1oMo3UoaaZM/0OfmaSaI8aea2H49nuOKblwHkYP
ykP8A27vmW3uxSCkx1kzYrpRpsiF5oWaF8KZJSuG5u/jwo9J0heSkqVohWba82jPdVLo+fMIs69a
ZBFxhBkqgwi+/mcL3va2JhZi+qfdT6FnMqerS/jdVnE0be3QAiGbm4MtX1VSqM5R1jVnLKV3FqKd
S9azN+sE6J5FEBV+OEAS1W6y/hUbPgsktw3RrWVJGwdCzrJstiNsVg6MIQuvGdFccTQL37QGqNsF
cHfkfGX9D4nnBH8ggbTXrWH2a/lQO6JEcmmiap1UvXVDBoRHYA77k9/3/ik5lOfAa1prgBNCokLa
gNLSBuN0kpS8DdK+bkAT0ah8g7SsJ9SF/4JGWeFT4rtk20BG+P/ZwVPYvEcU/mN7D+0wkTOiogVh
s/uGDfVu2fvzN0A7v7CKso22mP8QW8TqKp8kjetDow6JQrmYRFjrclrlQcBbLkZYk8PYPoXkNnRQ
W+sbc4VFAjZvzEaohfAB8ARNOMbrHld9PljVeXrw1AYIJMDEoRMwVlKgcZ70xVOAQtkHkZKAYVav
xfY5mmxRN6+mfFAUy9OZU6mIPDnfTOemVzTCiiVYyzu+QZoh2UNd6Ug6a418sxkcK29TmA9Y8HLs
UIjxaw/I8cW38VRq2UD7tqQ2AnrGuXfLosm/PpB0E2sxau2ci8laq+uXk9WEH2kgXNEkkNl7ZpmU
C+qx7mI7mCwrHnG44VpuDXMr8358uwGiuVew2Wd/UtsVDzNHWIdGohLGXRzfyjmrgNXOFlhRAkt1
keMik0xEqMkOUotirbMq/b/iZZU0Qs/dyxk0fp6sgP3u6S+bbsGwK7H4QowB9wIj6q4MlZFCIs4u
6YEehaVI67AGnn9OdGuztuLagSu4ffqi+KjaDL444pMzg6jpC8A3MJ26I5tOQBg2vxE06WxIM6xq
fK2jBHH9qdlrtSLmdwjNsdh150Pj05ETo32C5Slm3uUJDIgo3rDlhj5wZWl/Z3rcdxr8XSePBSqW
WF9NSuDNhAQwf342/3rZTiXlvYPOX9YpvwJjoKioP8gYXkMztiq9EDbVyuSqUOIR64qDq3ARsYfX
ETAaMIfS5mqncndisYMOkzGXYjW+3Twj3NM6XAMTmvOt3JltG2N/4uTJbFR3helCJf6CNuQ0Up5+
NGXceEvrfh0+X158TsS5ZpvAuGoRdgAVKu3I2oHnUWie6ZRTpa+yW6Qkf0RqKmhXOA5SC2QAG6Hv
fIlFNCsyFJj4Ec/qqbJF+/nPaJJ8Z5VCuLSr9nnQWH0qi9UPzWJT3X12d6Yl6Yje7ln2zjMrPmwE
AkP2Pp+jsYhKc9hm5KZsV7a/Jk8vKkIxy1pjghb9FTlA9mN7cvG3Xz5R/ev11knaTHgUsJKKhTZs
k7VrL0+j0JRHc6AbJjfCUYT8F01Zwq4uMv6ju0SyMjM9KTCSQWuTYaftziP8QqRFoq+XKmS0xFc3
L2FAK/PplPt0s49NJWmRODFNOdsPzAxbo94IrfkEm57HU2I93RmxNsAaxDYLgtz9tnM7oyN7m7yH
/LNzY2W1Byq+PizENTrUR8T+hOGEHX4CwN88mmE41qyb8vEAIfVOzwCBMJcsd4jsjBdfcO5yLAtL
Xm3hYTPprOrT6d+6yNnbki57t1j2dBU5sJQ5KrVBXhV84LXt35VlS3sEfAPd43PQP8yk0BEFaDzB
JXYLrlv/1wbuhJXLWZSXAxZGEPBh3pr6FsCcnX6LcKXfYvU0QS0qsAnq3GIEz8j9fEAr8jfXU/gJ
7m4cfWotpuowtU72mTD+1GaHeXROnANCsAtNFH/mdkl50wGqdf9OdhT/iJO0lWOX/mZ9+/4Nvnjo
67Hcnz9u/k9FCCIlV4IbZ/kLTA0NB+oUCPG7hQRQbgGnxjMs2CMZYiuNLo1BhsccHd8XcrJUE7VC
BFPy4moqWsc4p7TtkcYZeho0mhDasIipPWiUnUaKAFuwI808v1xfrWkqSggcJp2Ffiq7050we9Ki
7vlvGCSzOFmJWIMsx5hpRM4fuDCl4z8g0M9SC2HhVmCL/k0YeNL/cpQDtDEVIRIXZZmFQlP9X+1f
ljzmZcOItO+VHK0uCgRKXkaLHCg5I95QsNUNhfLcCu+xPBncxMyMagOJxNBBgIKJAw3YRUjyUaMe
7oadITL+W684Pm2kyi54tCNKnjZDHaAhBo+aaVc/RFRqaJlNvvc1kVezoCwYlqL0qz/AIwobWDMN
cIjl0jGx0sc6hAsYk1jX+FLsKwbiy1GwCzFHLb/XAlCG9OAq0t8cINXxrz/09i7eKb1BDwMe55+N
xUuTSFW6XF1bH9rhcJYo9Hw9AFZEIYWzWHqQQHW1G8oY3s/f2XKvtHoZkArO/wWNNZPYJIr49qEa
A1YvcYKLvm4VBAmOt3jVwlEXs8fO+QzzBHWqzUHWsxh6kMcbtvjs23zyu6aSPb/T7S1kT/DpHXGP
Ee1pGBpFEaGx5eS+7BO88EVf2zOUTQfC1X48KCgv4vwoherEdVCQVF3b0ncdgBrzMYyjviDavvj0
IwNbW8KSDsLFWM3OBQlL/ry2jlXvPkiJyFtV/rzxsUQO5Xf2RpUk4ZW8KdZXtkHM3Mnicey3Yb1e
d5Bef7TVw6KaOT6AXxz/J3GrJTh0oO7H2wlHbosFJ36Tlv+NHyHxJ1CSmPn5CqRyoci8D44CkWF9
ePB48m+UmnVtqFkpeLU1o+EG8IvHSS5u/wRlfW/2OdVfXpBa0GjoLSmHrDJoLMKIr4eUfLjxbLZG
85fSnTso9RktgCrgniN+2ICT9pI0eqK7aJJwA2PgyHac6ppnd3Vw491fvChLASPGW9iBgD7zGoSn
uIEYAgid19YxOBmAN5KHNfA3+kMACTPkUw13J5iArALSrQQ7rGedbAEVAR19BpKzR/GKe+1bBrU/
GLMss8DaqgLTrXD/ZYgMtfaD6bb64X2b/+bl8YfIT/35s5H+at6Fzn3c67EWToYlyxZL4+0qol55
UWzCWZg8yUODv/EYBBFr/9IqoXiGH74M/SJtg/Dx63TCrfPEel+R7ymrhm6mwvuI+P9TVA4ywEGH
Uw+3iXVdlmwZhDwieR98Abpk49AKvB4Nqh68aAz9/sutLE0+zp4YiFk5l+BGqRHnOlk8G9r6W8RU
0wLw9IdnhW53OH6+QrAlH6KqwMd7nuZGGDHE0KhMqJYkQymxs46ai2aoOLAAspJcyxKdKiMekpTU
44HhzZL6bWgjaj6iLrf0AOUU3JeU50dO3K+rE1ruzri8iqmJGtak2cm18PYOEVpy2Urpmd50kwpo
Plyz0EnM9ep/HzCGFd0GCHfy5f1fhcFPpdeQHTrr2pLonlFVxBBgcCUmbxA5bEtwkeafr11TPchO
k4WP8XA2QAcJufDy1t4c0mNgFooEbhnhErf0FKjxmKMunEAgqWT62a/zos5GSrOLTlSTACmS/Dws
AOVKJOnIwGa4WWcp9P8By92/f4GTPvs10TVm6Z9Xw/MmqBaIC14E6N3jGWoRSF20reRMsavya7s6
cFpQ6ZgD8dhsTIfnwwXCpQnBRwUiPUA8aagJomfYXvKcUUOVPSpmQQIsyhnKcPsy9t91e6RWN6ZL
ZrcYF7d4EC0NtzM0wZgczLM31GAQSesoG8pAl//5VALTKeF5pNDtpvcakizeEuKiJujmWyS8lRuY
rISNM6JtySpcnKNcfPMiNdz+tZe+DJeF/B+kKuMe7XAdPbGEG3c6ctLoITc51N1q6ioQG6fx70tq
37L7ZNDWDYUQ/LKFHCEel5u6nv4xUfOrZ+flW7wML5kPrV+XGofLzbnDAxRCDMVW7wvHXTnByH8G
z6lYed/IwRbjBgvGW3mxI3b8BEdBuzsFTexYrDAHdIUiJWUI9HNC5LO+ivJRt2YV56gnwEF9/PsU
JhNOv5eYCgd2lK2f04PsKC/b2SUkhL2tn0Og1k77v96aT0rRI/x8O7KsbtHr3tcLVkHo7d8w3d3l
p5yviO1rbOh51iTcMm6ACyjL+YMZD5fxwOcU5KEPQB8AaGQ1B+1EESQTjULyZC0Ub7HJa4IJb/lO
dm2c0Do25/PgBrRIpbXoQgyze7QwVjxJfy2wbKubHtXZD/nDgfZYKpiLqA5sPWde3ft1IXQx0h+k
Z85zb4nx35FZctBUbGCBGUvXa4beVH6eKHR42R/wXCuGHrmE1bdro39IC5Z+7WBP4qWtH9BYFLTE
9hRqHmAakBLHilyeMSPtqfg+IqbeT4EnL/d+64d55maEju4876tx8hKtgXmN88kg8lNybZI+aL9h
CzoYQOgrbq4d2K9hG5RPayG+G310AMVouUqanaupEI5DqI0xMPPYDFMe21ZuIoWFFwu75CStOlrh
1hkEbktODx/z1z2GsDWchCDFxN2bkeIdaDeq78+2LHn7FYNVjHIamQmkXDYJINHANX2gOMwDSpiD
0Qs69izXYBvF6g1ock6Pgtqh/a8zGuudPBFll1JdgPcVjI7/XNkJlE236XKRkcyiLgvxJm15Fhmw
VPLQ6B3ypH/x6ZcM50WYEllDjmpwzjHQb1SwvQx/R+GrCLT1bl+YTkvjZNMgIfGqjGqb/x6T7Cu+
JZZHIG89PPmEjKKOdkaLukKbqkihHhx4iHRy42LcrOssOZIyByMifkA1j+Q+Zjn2aaN9rNn4z2nS
RUQl8W+/M7emXzyxJ3aWNCbsNuJgpiR2eL/9X9RHBH1Qxw01PBw8BpOoepe9SByTPcOMkAVXO1ex
rpUjBqUSp1+GUCBd0YzI+alEzVF+8qa5L/kRWBRawo4/2MPs4d8+eYPRaYmAu248/eOS1sXvknpE
+toFY8lZh1V6YkSDpp17hEcusjTL+d8luVWNsbOs82zHe2LrfWE35eFPB4vveqfjNrbG7NqP13lF
4uVG87XaioP1+9+vT98q/Dh7xNczU0Wrje5INe1km4Z54iU3aqTWb/FDncPSaGCBY+QoYphN+WfR
WB0W3jPf4xW/GI3lsfrS0J1W9pQj0z+aBHDE7Bnc+u1iCv33EOsD8krneOl3x6YUSDiAuNPxCHFb
VmGhLHpreYoRejUza1tIOBGxIbKuJgJ4w5mLunFBu7LjAnYtMomfyjHDjTiXLeKQruI226rcJQkq
6mXcvdXIvp8ALq4zSwirFF4UrtYOAm2bk5CqhR3rBYxXvddmbe9OAIyf2kuXtbP49hsFVjHsnjXJ
AXyGYyi4/xFeDMgZNAudjcgkCwNdfk3szarQB1M5mCPJxpcSTKw7AjoeqYJX28PvksGpJ0BEGbYn
q/kuVLKJaEe4zFfn0y22Yo6VwaZnSYy3RQd5bDHqxVcPpFRZ4Bn+UjpPyOnohdDjuhWVk/gfJpff
6OeAXeFkcl4pRGT1FVJRbrmbjvD4GSX+JBIZvTzusZI5chd5YraZ+BHnqQPg9r49pM8v3UzWFbxE
E9qpOVn017Vwx8b7qvfeMsuO4cfl7Yf2w3vJCHZqH+2ImqrsJUCIcgp39hAUdRkVfm4G19ntugdX
oSdgwmTP7hn8rLZktCY54SOyO/Zi6q53hJwOMOOstu8d5SzKpTP8h6+wKVUwARuMZtrhmIE/9dxo
oghAfkT2blwKN8R6+k3uk7YD8kWqhe/XsWrqzlHiRaY80iV86ngFM1PCy5yxJy2n/TFF6KK4h5Lu
7O7GRFBhoe1pS27eXdaiNMkWN12zG8sE7X5se5ghyh9UEetjvTDrcLN+MeIUYUwtKQzjXRu/ZjH3
Mxa7Kn15M2OzpP9MCogO7oJNZ6rn7Vt2TsrVasAd0fdn4lkH/UVZmHkidquk8Zkm0xoIg6qNAL3N
eMHVVMVYCQxDt2Wf87viprAvedsz/Pn9YxjtDtRFc+ZKLSzdwlHSdtCDxhrHqW3T9GxO7/7AK/Zk
o4BoJXkkeyhz4IU7xXSi9OCJQnk/Ay1QoCS1ch1+Wbo50vo4mcgijTxpTQ9piucS4B9LKCL6PXE3
77jCL6bCvpIC1nSJ0e7kzOPMUdHxrPShUqj6ZfYoAb//SQWGsjaqsvzbpHluelBzurXPFEgupePw
m/4u9ewgjg3MIucoictGMirlBLKn0sLxG1oNeIh6O/d785bDvRkAfFKtb687keJ8DCv45dfj4NLv
AvfWh1YAQQk+oz62bxQ2a+vQ1xIqwnPkgC+nIc8720ZljHjK5aZzmsQhROlLr8g27dHFhX8B94xE
wqDWoBTD/1jgPnxfIXn5qzV+xJdUw0qALn8nml/82q7X34Cg/RVsOmwJXalw6/Ihcpk8k4Fh1vwh
5Fq5fqYpIfaqrk27CJmWkDtK+mZEKZUSiZe9JlCMqd0BE7G4qPAYyCsbRE4MnPFx9LbiT1TJWNku
zQKmKXhHoFJifT4bpNF1uVYTyvt/yMAt3rihgNneg/SjFmWqC0f17jBiWWsCnSet4Mnle9ZaJgPx
IYz3bVgK17QmvgRpPUDYFmXpesi+NbGkrpUCzvauT452cNfRz3JDB/Q2k0hlDqy9+qOqGmpzz4kk
W7EOT/M29xADYUb4/Ml8wMsxpwP8rTYro/cYchC003tTii6FxcApiwfrHUlvGgaNHsCpbs6HpclP
nlBBVq6AunVeTeeJBzh1BJbb3XxfsFqYQba1HKJds+iTB1O6EkMWJTl67N+Ka0FMeO0Rv3XNE6pw
cko4ZOpx65GVzIFMQ27XVpTkirYDn0QFdOkGyY+aUL2uWh1+bH4OC0oAmOLZVwu46+mFat7PJPr6
insbn8TRM9S7AC9h4BD+hCoWmr8XKQRkvoaM6WPTqBd1JGaj53myPfzGSgWsQtDZZhgj5xTv8Kg9
5Sb4KgR6VED+PFroKMmVQHt9KckIVWFx56orhY7AINBsxbNTGMrNcl9VzwhZHaNQQzvMHKGOE6ww
eISyD9yu4duu8ftq88SUMBthsGWu3sFHL2CXtDtfX7fLM2qxix6uCEzE87mu480SsdUonGnMBJT2
5SkmJMEZxIvbFM5Sx6up2avYgWF+iLN+MVA7OipCt5gJMdcLh2dwTfFPyJUiMUZp7B7qnsLIZ8tE
hGid1zwHr7a2yCNPnc68+qtB03TBOauOW/5dIuTDBOg5W0pPULUx8pXOIBEDRzOvWfGppP5xvtw8
mbjO8l+vU9SR1hL9zzA1EQ8KVk3dCpNU3bJoIgsXCjIsTU3VcLtVyFYGrzKpkGGN9HGFStbM2fX/
O+PIp9+I1QzsVERWy8/5XPU2K3n0OqYfPhA8Mq8BTUIl1gSMXUcudxSGhwxhaR+4De7o8BpbYXGf
SyMqMOm+TEjkntx0yPrVrln1sCidKnnjrX0apVj3YboRyVmIVaUurJ85ICS8OPCYGXKDauLO7v+5
LxEBzhfA0UZwiJh1VMYbYG5zgNPXE5hpTda3VZEDLgJdP6pBiWL9toW3kOMkaUtXdxFeCFPH/iyy
E2t6Ureklf0AFxNHlu5wnIHYXcvYtfseCztGc1VPtkAqbACN+qN39MgXxFrEV5w3G96+r1Ox1BXW
gwf5Y1v4pWaVEduoyyl8GRsg/Af7miCinGj7SaPSO3jdxFTPsVEBmgKylpFaYL8PZkjsDiwS+WQU
PEvnwqeZaUtoMBq/YPjRS8gqE9YDrO3KE/8XzSqm+RyDpHkczSfTc5dyPrNx/LX5x3I9nt+EBz9E
9zYt5bI+9J+xGvqe//EKbJi9kU86eTE50Ycq4zsKpj6kfTz1VSbKk3Lge2WftW0ix65ZbhqdbVgB
8XHa6qY4o/eohdzc+SDOVHVTTU9+5tq7mkRZCrGBC+SrJaorx2vrkd/4Gr0BKdKX0Zcj5jUCL3O5
//YvfhGt8+9PxI2+4SbSfwsbvs8ulvo5q6cU54WH3mzG5Dn43RqVfqhrwYvk+rGp3aGJ1eVxx5R6
7RqaEbjcfNrIznZB+pRkMmM8qes7Uu7DIjLm+Yfxuq6S1EeznittHgQ/GnyILTLqPK/+VZh89ic6
2HqLLSA75HYculHnRW50Z6xVYXZNCi8rYTqsCYRAGGE/5YMKu5mvzkknKIQzJKpfSGQhYk0u6X/2
LifJf8/kg/mLSi9vRE/s065Vn86fzeo16LbEspjsgljOkCnemvwKRyf8Wn7b6aZabknfF7oITZmj
2VU0Ag85y9a95S8PbyIJhpJliUtD3y4OzHCFqVNTozwdD38osLfIKWSuDfhexzKVUoj26oFNvos7
3K2d5263EC1dLGVor90MYRMVbszoN0Mk2rajwhieebjm0+f02RS8u4JgTlGf7ZQvQ3U/GQF23YTz
fk3yVVJndLz+ksAWISTZ7JXhWdd41cvxoOEfYptvqViGnj1iMC4AZ2Y75ExlfYsA3iUiKusE8ri5
LygSTU/npGZhls/SqJfxb7UYexvGsVOlt9ObVHsZSIUfJ23O6M2QvZh7cyvZsxe1obdAIBu57a2C
PbIlRDPalUu0Khx8RvLCp1lieu48XK9TelS081AwBV26sLdv3r0LT2QDL5xNH9jvKP+t9q7cSVb/
ku2QfZVg50aVmeu6fqfxYKR1wVrsJlwteuBcdPBr4Bo4pU2UNKGPyFZPblYXe7CCSCh9D/44ea8N
6zR7iRdMZe/r9ASRA+o8WJPS+Yg5wrk7pRLcMxT+D8sdeRNhDj9drlZH+mJ141nCEmtSnQHYqMY2
TK+VHEmSEWvd3rXXIHiJIvcyYqMQBH8V5iC6wslQ5K9GnfAFEhtG03SzVMH3E70JqKW/UFDeKSUh
rMeUtGnouS9PwsLyPGFdvaY9AAM9WJgtFu9MO722eNu5sGKx4ZVnnpvt/mfMwxPHWXxeR9iVWz8j
hdUmcAXau7DS4y3R/CGyfQ0I4w9h+BdD1N6J8sMElrpil7/KcRmloviLpU0aO4Ih2gCe3pmLlgnf
Ju/dphNf7Ejivyclh7ptpcCqogSLh0cmrjU79wBDd9zgAIy9omA9Nv3bpFBK9ebmIK9TMe0O0WDa
zP9ELbppq8GReCGuSdUOS32O2yxiym4FZeyJMLykRvHNlv/OaFnAOT+luqay+dOSKIWu/roJHFbb
dJAH2UORv0qDDKaH1Vb/XtTmFIiU43VtZljY9/YI2olnN6ELQdnsW/rpgMY2xBRo95fESsHBl5JL
AypUxtqJV8PQ7RTmgSBaxaXnpOfqKUVcRZzgdL3xotL1ISC0xETbtBpOFaifS2tNV2qjWqbdEj+M
qDf4zTf267CaNt+cd/dD+oGzmaLguIVMZqMd0qbUSbF3cdJ93l5XiOstgZP9CudB0raFPcQwPtLc
Sy5McDRlPngobxqH+77W0lSMRFRSDQhaAhfSidqUICXz5E9PzFqo89ECXRhVm7NlQZRIXLATqTGW
yiTJE+M/TrwV2GhIS2ulzs4kCDRibbHPX4OoUC6L1BFiCZV4Q6vuXtVmKoZbVP6Xjic19MEjs86j
7eMM2Nk4t1bOeslq3UXXppOuGsFZ8JZ/0/20krpi1aqwB5PMIRxEyRrvsN4wSBf00IO6V1gsJd/m
kwYO0bCSB18SeJiTybTP46e5WEgZBmu/r54dPruiC064TOx5KB0cIPXNSVfcEEIxxHioHnNq2trg
eawSdQVwSODt7t4ouBXGhAXvovKTcIsh0tvveWZzm0/5Vg+Vqm+d9Ni4SLjZ8U6DO/3EQPhhSo9S
X+LIgVeJZGOfwmo/iS/rgKkiwUQqfTg7PP7191wLMK9hrTjEPOAT200ac3V/BwAj5fEosJo8FjW7
db33J+RjBAOS4rzS/SuO6xcyLje8wmEBhcxBnLyS6OGyYqrK2XxjmAQDl9DIdHFPUJRF/NoUv/Kx
fI9BrLshZ7n6UoDerQIeL/g22donPUMkZRqJ7t9PtpHXs2r462T6PTl06lo0UDV1sWs+PHYyffq9
WvXQKF7I/lU+o7QlbcerSDYOpDYqq2ySIbJhwQ9qqQRke1w+VunFx0Z58ipWzqlrgCTinu3kGZR7
USVVpbHdXPAMYe9hjuNo8IXEDJJeLg6wRylo0hF5J9PkGB9I8p92lmtJd9t/pTvrQXClq0+dThw0
LSjLSUogPSOaRNHhUeKsaXOl3QjE19mHx0MbYZQdTvh7hnQ//dpxmpCA2NQ/rusMPLxeS9K882xE
rJm5vpRa/jLGVYBJbA8L4FrQ+nVkkSG+CaliO2sgPnUaNT+/wLJzb3Y8EdanBO8/BWI9T5mWSxFl
8SDDIj40BSOs5ZHutfFCF9eq8kGwxgRB04aaYzIlZ9QIU3rSW3qqKj3D8B4znNwEdxbKfgABhQE8
5Iml3xqem1lYrype0PR4r/ya0f28tDZplLZPR/M5JDoT+isN95SZrfEWvAo1BEBSmvCIYCorQFH7
5mWdOFlbHmiokSVZ/kN0USV6u2m+d1kO6/u8muXyrNSAVAqu2609POxR71ULLwlIi2aCVZT4kf0b
Jyf+b2mlXlzUnQjGqPlchIQ005ThXgXpLoNiTNSgGcNfw9kvfJhCRIeaIO0zDI+oJ732ohY/LE8D
ofiCRKmgDOInJ7AWcQ2dSe87ZMlrXuMhhagTI899ADyJrNzNI3vS2OFYfz+oxJFyOquVL691h/J3
HuCvhXB3MSmMKUk9avBK4f0mzKmfux/P422rxRR52rMiH9rwtXWjw+uBHmSCbsgJVcVMZi0Q8SvW
gVGI/diss+1WwoKaCcJ9feT6DyVZFAAtwyOig7LQIUThsOY1v2DWBUEa6IGxu8grYVWwy+4FWbPr
kn/EPXDWp1wYjXX0dPXuCY/mwqiCtD+3GzbKgZTe19Tjl5/KfqIsHIREMt1ZcdQqXwIBFyxZ3CKB
fTAo+K4mg/keipTo7Yu0YzqKavDygs+zUSROTYSt84xYFoc9OLJBtDz2fUG9647hHoRDgEOB/i0Y
E8aFpyvVg8RYIG+imxHCyY3sORL6g1DnZgJ8DB/jZz6Z21bLxUGSYnqG9HSDe+LnIQZj5b/aRVV7
AL8uvovID/g5CAhEYbPeEYYlGJWQKXkECSsX+dS4nmfc2IRUcSYPmLh9vGeeO1jQSg9zT5zUSiKw
3TgeT70oBPL8sh1FXsHsbCqFA9gGanL6TEyuU6BScOSB0JAqH3pw6MBRULioF3UtLp+smCAzNk/Q
p49WJoJkEKs/WYSmKwCD4gXoj1vJ83ZYauctiyr9XUWXpVjP6JWlCbBoKkofpvJ9TYUkU6hbS8LJ
y0nc6w2fAeh/TL+gvdykvKT2Euge7aEXduJxhwfM5uGe1WWLsoYystDA9UNcgrSPAqTqtsKh7nBy
POOLx/5ktfwXuOx7Wp1GqgXpv4CHtmBP0FstDuxq9rRA5VPrSdJQLAKFnxfPpIAsBmcKzuuhfohY
ZYd/3Qjkp3gysX8iD0hZmzb8wv5zl6djaBVgZMmwExYqcv8bpLzZ3oIQ1xbEfTcirgT/uOLWI0Na
AA6WXw8leuFs1l/Z13GP0b6d6C3yWTdUWkkgVyzNttpEKSdyo1znKhxaZWppS1W2F0dpuxcavLqA
5lSAoOtr4H0HsibwO35KA1g6Hhjg/4emz1txdASiJ0IoKXkKUDJqeDz2BPYtpLkUT86Kdj9Ooey9
SHAVXwasuctV/pqSIiWfVycSHg+LAQM47Ubzs9ixgkHt10ocw8TuIk4t5PdapkIwO6ZCdWrMAocp
OGuY/N8EqLDrlJoBokUGeycfmzYSCcNM7t5pR8zYktxhoZA+OQclxhDs3BTe4WALqXVjdwM2azPc
EJ/PW/QJjE/CITRiKAE/FzUzlYUAUFjY5cvL3R0J0gVdbQC9fMOxfCBnvLe+azswRDYDhgwDd7l1
HYdGqW5SlAoPii6OREy0skbBuV9PqquI8W4K+h2jSPYFBW33G0SW527oZ950j1mlknKxCOpQbiTY
gfKAHWfFS4MRuolD37KnxLuFfxk1EPUlUPp/u1VzDjsvo3tZLG3POFjoBFhvJNNXD/fQL3981Vcm
ELMGU3Kk5ESSdT09gIH9Aa4mW4lQLSeywMoKEjWjquwS3J7xstmlyw0PJFccsStCLmyM5lT07/4G
3homDuaoErSBSPGYgd/+F14J8jV/gC6++iThm//3pXO1WHzZ/gt0qd9bWQsKbic0Hr34uS1CEVa5
j1EHasWozb2RPODLrcSjsjr1DbSEEJDR/urGMiboErSEx0tBWk7ynLmYxcAWxiGeGo3xIv5UiRoc
ViaF0eqAouPKlAq50nUtCkIDEXNWo6Xn84g/pbjuq4J7h73SPGDzbH76Ea9W3PeWbIi2hi+k8Ym1
GTGViUuPUDfJNb9DsLNVZxqk/+8Iv9P/UyMg/OKUW0xe5x3ogF+kce+JPdELFtKadShPe8dnGEUd
9FVW8gJr4BnaxfOJR+RBl1FhEOllrKYYmc+5FjbPQYb7+Nx1RGdvGkn47ch94KadlF9a5OrxROPO
gKBYrOypwH3TvgnEvkk2HA90IdHxlLSXnksBFrHQOYUgjguLT6su5fXMUtiNkuNZJLe3xBulbLw0
zzyLd/HPoOd98CMF5Bw7LBbgEmORL8wlmtaOtlF5DpSiFdzxp5cywKhDiasFKZnk9oA7+uy/kTan
L8tp943Gbrig6w36I5nCW2qjChnX6oEMhrQ/wSO0TkvBD+micXOZ7Z3TmlpCU6RmFaK1fe/qSWmY
ViZBDF8yT8xKeVnGEKpfU+1IDuaUQmL0yRX3M8ggLf6z7C6eHNHDAiyRUuoGFgCKgmjTG8aT7oOV
xK5Kvh37slO4M2FwoF2oGQVpcV6nRvtnC+wrks8sX2kjHL3yF0ekJsNLYiMm+mr79KDWYO/CKapS
BtUlIQwGsp75vocHviEDEgwiKQz0krgviBdMyLSQ1IRRd25nsit5e4LsZu8DqLuIEjEznDoAb7Fc
irdwdCvINEaTdIXZZQPCarzN/eTbN5tjHTg+od0I06B31cA4Pdjk51jJzt/ytJ1BcJjeCRNnAqH9
jyKPLa6+3Hs5LM+jai98VTftMCQv+fZ8tx6F2r2kdEIW6+Wb3WoEwpC/QofkVyW3q+FT0JYwronr
XIZ2A6mB518uL9v8TOG96mvIzfegnGznn+aZs7/M4TV5FYreOXgOfLomokqLcKLYFIbPs4mxsjRZ
UTBoecx+WujHg0F5C/wDGfmWgfQ7tiGo5gfXGdl0MghNTQgr5/+Z6u9ZW+C0BOlYBIfZzDlfLyQ1
dCusTrLyyjksbAL4dpeOr6zlkt1B/zfNmKnJkMbsRZmtfmLDGnarnRs2VBBTnrcB24CZR/Kc2C51
qjlWa7l6N2Y2hh36y8gwfVu8kZ35+in7f1OC4RlWamykxi0NUJYxGeIX4MOv9QYXK5fmp9BY+LLx
YjXb1jxBcV9QCbYd1kReyOUYMd2MWbEy1grYADh9+dpyzwtsrHvYzNnVFEnB7KMA3KTqyMYnT6Q4
DHeJ//LIlHMbzMYZJwAu5xzWR1gvEL1+rLNx6pvPddbcwwHqD8Z/dtzu8iZkb1eIKOniunHP30gt
xYcpXbYc8ZTrBSDEWpdy5mnQ4v3XwDcRZaJQvOsael8XtMHoCLtfgCgznqPq+QRBxkDlbOEps78B
m5t3ABtJtEhNSsMjg5WNeWCDT+d2ee1lfYueB09TUKCSg6wgkSIrIOxbQYNOIxlS40ya5qCs/c2T
xxjoueAV33YqGtcc4SWTSZ9xq5fYo2OuXbTzq1sW5LWumwM3VNURaV7lGbs5Dv3oDpOM//vWYouO
S0mswHepFyfsuENNjJ/A5Zlk56NC0zHZFRusVqWS2XpoCTLf6g4rHzV7X1b6cnlZjlLcNAwhmMdZ
QVlkT67W4MxvQNPOl0EprOXiup0s+Ewt7u+RGY+Y+wM0JuyoWkfkn4fMgpI7dgTEfL8+5FOEqspD
HdC8ZcNMaYTIRxn4CKhOgvlB4CnYluL14NgeQXK6Hvbvs8ImIbxCAOnq60bxLAt04YiSNLaJuTNz
m9vx7sYpl5Xy2pnSwDfAo/+TVRLnrL5osIg47v6WK/KAOwed7nLvEoG/WpfLOk7SbGAizxLjjZAE
33+A4MdsdSiIQRZORi3q0rsOQjYi+bStwM2Xwf8u1d/4yWYAuTkzDBkekyCoU3OYetaLhqrYU40c
zVFYaTOatKqfZV+BenjdRQ00USBpLggUNAPqWVY60D+vvfqx81NlImwdCtrMU9/L+2WCzl5RexfM
r882slaz9EUp6XN2DBHaaqKtQuwWeqQjzfIoMvZoHYHmAH+YDsfTZiAi0v6/UBE9svNk/XjzNKdU
tLre8JccFi27qvEZ/ctzybfeJWlQ4Rn+nZr5z7wM58ZGZzXvoBtp2eNitKtBY0Fxao/Ps4lg9wnX
wj0mHA5BHC1XOc0HyMF6YG9nuN5nhXg4ehrxr+7SOB7l50eg3P/Mtqc/2lKIwxlnEE8N/WFN1T6A
TI4/ZR4FgA7nMq7jTew4LaJ1TfkhRjmViu6u+SZY6AArAt8nMzdh+cfAx+gz80hwwpbtgyAjJxzS
peTtZaeg2zrlQU4p3n0ypjnpnjbV81EKgSQTrJ0dCE600OR66vIKg/H+UV+HtlBfDdIzC8bcdLSt
NRXynTu/EkmF22vDW/8MzHPZu6t+jlDoPMJaXk9uAnGCJFZmsr+IH3CGbPHGCcr8FO5sc/KWXk94
XjXz8hyFNOI2g7Fhj93toJZ7UOvF46oU2eZcWTfBlTXX3X6NsLJ0jZxZUPiHR2okDQWsZaJ1O8/o
/003CJVA1zugbdskGtSBV2ptWyrcUGLGyakUD8octM6QbRfWJn0tDyrUakEOacxxSUkB4lkjwhsb
nelPvb6+4KW83TLUn67kD5MrOjqRoCSxYtFvGTzD/H6+RGmqGbudn+Cc1zUX31zdcgiKBpVmRHuz
aiy7PLV3PFQ8zhMUnAnmhOCnCP5+fIhBY1nj2JzeAV+ZAHcNkCvavo30qdjoKwzPWcpL40GYQxBH
rSQdTBlLhefdxhGUM4Hxb+iKBbNJ6at4q1cZ2LSni/bDAN2iZFwlqPFEoEaSbnPUnYQKTCMRJ5uc
SFFQOVLgcDylwtBuVXMv5y7m/NVAe+XOd+JKwbKBGx8U0D0HQUEDD1e1coQMCwW5Zv4hJF/Gj8zd
/2IZGn0EInjZhjJTjQKfyQjpteuX145bU3nkch2XxmpUH4ynFKtlhEsCOaAaAn+3hcSDg9mUmY1v
wUuwv4nIAuhH99tt+hL5PfH1p5NKHjbYTovTlXVEFU7tEFTdwUnDGgkKLtJqPT3uhvFwIjWkj3U5
Qpuk4+nagRB9QLwqxUgGlXcAJR9oEEIjjqzmemoxNWMaCNTdmdNrjOBTzCO/xJZzCGhcrMwJ/eRc
04nHr9W37Uc4Q4vDpWqbk2WCa6tbxzxtUlZdPZf1GlSNfWqRM60gNgbwF4vdnA56MVJQEL7Em4Bm
0w7fSVriEnx+eGldhj9/j5Aj+PuEVirawxWZe4OLIqQibxn+aO/mkZN88AIkwt3No20HafLh28Uz
+PFEZs3YPX82IYmGZ6skMMyxdv9YsMf2As+F3j+b++Jbr9kITcNYWEACNHUBhFYGbbHpGwiSHfxy
G5oPGZY9YuvU4YAnpj8MRweMjVQA47S/yHTJUWU8N5l0LllRHbRUG0SznWKatMaCCyVYvsF77T5A
xOfetvSJb+UlmZh2GGLmc3bfjt2ycIiktp+oD6NRDsYloNkSQFqzoaN5YmZcDKozJThahBDeBaRB
VWt2sdendJxN97iLcMaUAo0Ks/3WhZje/Xa2Iv+QZH4cpUYif5mMeNJjGM5Dn6u94CrRQn7rFcqe
X0vqC4Nan3F4pZqkOs3P3F+hLeBE+6hS8vPEer4bGOBiVa0GeDohfB6wJcSfPj5v/B6p5SDP8oiT
rzmzw3Idr7VBZq+b9Jopu/xsNBQHKeuB5cc9O/yGYIhNKkkLlu0RMlANUxAYl4KZJza3NaU0HCLL
+B2uqaWSLzyrrfZ51Ugv+5yZpSfpejW+oYqQtAFfDrYqeEL2/djyoCnISm0SO17Zab46GGXhD63M
7h266vpoxrnHlAXWPRCz0/BFBgGao8SHS2mayIn52vmh8lVMUCMvxQTMDppApJwHOJim6yJK/j9R
dJpDkkigACSRKU7+mvO3jXiPTt34LmMGQHgHf0GlBlnxPVVogmd8p4Edpvv6yh8kXElvTJYXVp7v
jUrtF204dbI5RDOG0tcYnJX7IMGbMZQJhqXdvILu+CO93ElfhKFhdJ3M7eNf8oPsyNcTQAe7rP+e
wpeKBwSBsxcbtg2bV2IyY7UDLo1fmyqmHuDIA6zv792wPx+xu5t9CYUHKnbQ2bu6pdbu2fLZw2B5
fAaqDKvdse+bST+M8nAgpMbP92oARYXO1WLltpDAXSLHTvB4u/VkuAEbn9jV4sk/spQDUFh/PlTT
DeW+jQOemngwJ2hEceM8sIZeJOiRRlVXoXmAaQAdgclga7F9R3NfJC4jtusSQGxAmKYgt+1W3SUh
IvmyIrro1/kmbbpo1WNShJLKtp04q8A2CQBOPddX10r2MR82v77O8C3+XfEZHp2SUqYEPMWkUH3+
dLGEz+AB7oZk//dEbytT01rOZP5CKM/m3OKCI9mbnzEYiY1SdUVWSC9DDruJsTHpL47PcbfKWmxs
eQBF5XRl9PqdZdmirtD0fUPH2dHTG1/5t6shysKBzUeJFMw0V2YlCtPJorClBEprs/b0ZN3goGwA
rsi5SZRUim+kTKc4GZIFawwUG3ywmQyoHD9sbsExje/xB5Hc0bEohMlMPSOLcc2qNT9uBWhYs54X
Cj5naH1xF1GzE2Kp/qiJFPLdmty2rkWabii+fAKsdmvU8EUIIUmXBl7KoDxN9NWciXpSwv8OYqXA
5Vi8saPbmV5e2LJAU9uFJ/7XWwwy/S7DbS0UElg0A2ekoSx4EtzuStu0dkcyC4FpQniGH6qdjO43
ZczdqTKJxkiAoakLVDGQuA4CDuaTYB+wzjObIxozF4y1VZSpPMlJJSiy5gmofQuI5Brj9fiZ5qUv
28kMLW8xbp4Fdyp8x8LQsMUFmk9LMGmN5nqYegHyzqDhmETP5zmif92T+9efsXcbRqBZyATB362b
7g7I4iM9bFqmXUtSUyJNH8SSfZx+Ydu2I8AwGWWd2K1VFnDZarJptjB28SiGC10MrK8Fcyu8PO0G
gbMkicbTCn7ebF2O+W4qUCsv6Sv+LAVPepPrxJ8BuCnJjj5UPQ8TPE60Kls+0mSBUTcgZM0Kq8m6
rv2kTpGwCtQ2h4+jH32oozUev9YZwuMnvAGxTpNt3QWyOJsgoLpMpv6PzQ3De5KIMQ1ESxUgss/t
8NL1LehonGd+cTW2LAgUiy1gdECXdFTCdoMcoKzy9vNxw2U0ymayG35SPLkW7CA5q/y64LT4ppWz
jd7rJw3IuRVrRGwoBzmnGfpbuiTlvF3DU4ZzfDlgjqtc2sKIJySlc2wVafF/6APFu/FP5VSeUiQp
5nQyei3LB4DiQEbxNSan8O+dpmnbYnP0eR67M/KJnbVOwnd+2SVKK0qf7Op9kbT3LfVZ4GB2TkRk
o6ar3p0LRRvYfgSxYblM5Ezgc9588c3nq/BQMpAw5Wff4u91aFAhY1pJME0Xv57+2E5gbsZcfyzq
OGEtMqUAdpKAw5vvZ7bBkiiJTh6kEKBELK68jcLQArUWzNVB/VK/qsJuOOOpTeWvAC0lIzuZiXXs
MYCL4z7KpQJzBvHrLwvgdg+gbTxZp8cBPA1M5nUm7LxkDdtTUgJdxeCp/s104jBaT0qzv41ucf2B
JiEotiqtM86BB61cFLAKHGLNpu0ioxXFhcvKAW7W9Hen8Cf95uYDEWI2C5XwkZ1uH4qJRgfm9mF9
cCx1aQNKNi2Qjp7NBwrPrE1sCFsmO1Jy9Mds7Ad00BUuXDLPmOgIbQ8yPP/Nx7dcws6toy4iyXSM
OtxP1aHVhG34Rl2fq2/9oxLRuFxesFb5gkIQ1T0d2mU/V7e9SKq3cV27ZzS6BQgIhNBK571NlGhf
AMslugrGZC63tLX39EkouhBOErsVs4dMr0pmlv7X2yExcH5Iq/HUF56wl+7/D585WatPg3doVsRT
5o/eTPQsviKKVXZwUsYSkmE8si9Y+DQGy9B4qRc+BJuaENVTxI6VndwQR8xi5XjKN5eAaXp+xUIk
s5zYZbNAPy1ORxWUx5tNxx8kvDLNFuH9yhkUVivTCpYks+0GolYR+OqSkbBC97vwQS90Oefb/acC
1UG6dj0uGnwxS5h0r7VBsU3L7GIM9N++ZuHDTVGImO8K7yyaU9DGfcOnbDHLvsYDph7zJj0pR4c8
3mNk76IsB4Eub5qpxP8a7rHAc6z4O04BTsRD6tSNT5Y0XjunOmGIHE5k51oS/M86al9yzIFP8DvQ
HCaq5dLXjAHYgnM8SfgVclFKpZjXBaBdphYWyeRv1vGJYAKK1PG42mTh5KGhl9k0GztJTpZ6EIu5
UTEv+1shjqgYWLFFq3zjGnHqnJkUtmrZ7Mgg7cVSZ/IHlDiDyln4PVG4luKGjz8bEc7oDnGeu6En
0W280oYo/oMs8lfbNrY8kINJ7gWhfV4N37DqQWEAODA+mBUrDkBcyUVx3ZGjh8xrVdUSdpXF8HWl
PX4mqetlkmGjsiUyYlS0LTe6UyO7TKmEBTjSGEOhUF/8NoNy5L8UfR+Q8iTs117CV9oVbS2WjXge
O5SQu9oKePnpAlaaewB7P+Q5WQybOlRrFo4BKCyb9CVC27nLPpnLZV2BB3DwIqa66kY16RGGunp/
pCJGHYoz27Jeiy2BlZLG2MoYmUTQLpJthEw5KSAKyxa28atv44fdSkR4Ep4iAkzLwjKrmfSMhdPa
HSxCO9AlNEyy1Lkp3UDCntyPvPpv1vKSbYQDDPFvhzF2SYdOz3xqmuENpPcKndkXtVqYpmRr8X27
zSm+Ug0T2yjBsJdndP2/kmI4kwnXZky+fHmjCiTbLrZOKNLS/aQvhNpmCt0lZHXoZu/k3KR94QFU
Gw1QqoIxk0K59Bh7nGEONi1AwBhqYnwDvsVHvombFWry7GivigH+bUG9Yxf3tSqyeafLVGuiTgqo
qmS5zX5EZdeReK8zR5vQ8f83tvXgKWxTA4N7wA2bNQwJeJ9G5uHpCMX3Y+xdwP2gOR8AxscetRoF
3l9BDg+MUuBKnfjIxtC1icDYm2J5Fn2tVnk0lNia59jsXMPkUDMqnKkqPWnQOqJjJLvndAAXJuH9
aye0paceJsbIukcNPRiVEUPLFqqTYGohfhwEi7o97opreLXc99+tSXeYXM/G+0WyhC0Te3zbfAgQ
PZF69mWzZxlwwOSVrJPRHDUuDcIrHoSnqAjSfZ9+wFnyRvIB7nb+8/4lMToTc/c4fp1qOKzFMwn3
y3B84sjnX4l1HIFK2kvszQdjX0xZ7szwpZwneYDvNfNArViN0hzekR2u2Igpei94tiItdzrAtn1K
Fdu3h+4HJLZpEPB4DVX/1brSH0CQlGSrqYjsHLVUwLjcIIScu1QS2IkwGQ2ONxxRVQNIpw8Ft8ZM
0C7iBhdb4loH86LmSmXFclZiC/BmvS0Y5iD79rLidGnbdhdkX4+aI88oFOha0yS+7NsiwsAygJsS
t6bHcz+YmhR7L7PY4SjCFlRDXuYeY8j6U/Dwre5BPnEdLa9AuPHhS3EpdWxJksVDfpkai00FZm22
nTeWSxt1xtppaDfF39zV6Wtkx0Gu+cLnlIvXdfkOy6wcpT7FGtmMFJOAxeGlaTBNs92WUtFqj7z0
m/XBCdrfyPk2o6mBQCEoJLe8Z+CaH5bPnOBSsafkeIG/kQDadU1c9N5w80n4coGluhoujaykJHZD
5yzVZ/M4YB9HhdgB5dMY0lv6+uzIezJHfE5aEfeLUFyznO/q5Itzq6NH2Bc8ST0vZbBbQ/UfKyHi
yUVR5WRDycH9pyoYMkBUn0rxpZRINbfZg/8F4OP6TObDce8Ivo6mTS+Tg9+q+u42TThoo52qs8Hy
4bi9ZmIBJD13F2QVfkSORhTsBOPMbM0zrW0TojkV/SaURRIWjFdO2+xu8bvI8XM+M2Gned/6LDvT
6WosSlEh2aDXk3aoH+E/h69sGyWZRZ0bD0DXx53OGrufwLf+TLPpLW57vQpV/bvK+nghng5qoX41
7OwMjuX7FyK8R1qlIB/Ssne0BvL6a8kZdIw4JyY0JGK1LtXP/wuCHOcdeiqGRJ3IV0drCtQVwNLa
ijfT1PBhlRoGCXQ8HGzu50v3U3M9jdvqZvUTaeRhHF3IFT7T6kNisum7Qql/p+V1J0JR3HXEp4LL
Xqgva+vnitv1QX3uIL+JbT2wqlUbqEr9b+1iHyoTbulDe0oi7tncaOvQUdXspC9qHTt/NNfHzLek
hAPF0JiH6JOVa08Ct07qGBg9DgM9Te52UcjBlEF+3Y8ZHpLLy+Y2SrhTDqgdEJNxVkK+b+EJSab/
H9mWjkhJo2T9Nb3Ch4UOZhPnDavTmErhIPugOxLc9wxPn7KKarHSbGnP+IIJfdT5Ayk7iU7rPKae
ZKbwtOpTCoOOWhkOWg51ToiS76jVQErWXGJH/5P63Xnf90Vb+RpK/MG2nTRV7Q5L6U/NTd0I3+hO
MxbYG7D8C77/k/Hcl1K3i+CitKbns1WV9JEjH7joyzy8t8nnTAApFxm6Ez5D6wrVNoizvVhzK26m
Ht4hJ2kS1yO7Q2+1ylhxtLYU5K02MEMGvfq3aLFwQjUxd9Sg7vQEVG1a+BCxTq+l+8BUdSWANn9N
YCoqso5lZlBtTHFnZ2a+7o1hIDPx11+a8z1XH/ITJyktoQlnhhtVxgxMP1lL/qqOnWq6wZEAmFHg
GSahTZeaSuWRzbWM0K/4y5WMpOpT8yaLjq13cTDGNHKr4NrNgHnkq0ryxWapwVPYPAdml9bF9dVV
NYUrghBHOU4wVPAZXKxWe0glvtKVfUygbEjuizlQkekwyoEgxaawvlAiVQPK0esGByj6rBzjTC+A
6DiZRO1cSUaN4NLzrwHPy82l2C87ipFDQ7nEBSH+UrL6XyrBF40Io2oly48LkVrvWBP9HxXBT2mb
ha+HwUbeplqahYT4EVYaS3mPTv8YhFYlY9mBuE9BaXAcx0OJ/VOxrctRAK3MnUnrd+bFHiCyLf70
q4EW+LIZo+EIZeb37in5+hp4QcwMoeapez6U8Vx0Q4YUbKJbJ+joG9xFBKIkWtmD+YqavmXBSgFs
X7y7zHl0XAtgnnlD/hIqhIuDKJzXEFbu85G7k5myEuBUJDmlc5w8gkpEL9pEFNxQ5BsYbKOusMk8
bQU0CawtaDV/cbLDuz/BSXdsoDZjvrqtfNHknSSfn3/uT9RLlTsXuV72NJjpAjFv9ZkIfPiokDdu
QFmxXaqJ6X8nHLx6quIBV8ut8BlMSF2XGHB2dHrpbuf02ji5bbOU3HJzwOIjwKGernoa3JcsNPzZ
lLZwGcLtSYwcg0CkWqRqwcPAdvlR7PfdLr03zcU2wRu4KGO2FheeTYfthoLHDx++e+PEircJyfnY
QjmbA+rPW3ju5epSZxEaW7UeNguCOXlg8A6RCyA9iLoZ8jPIKhiEzt0qgTR29qUd3D814OUVgQbg
B5IBEkB2EiVvhz0SR5wwXaCf/lg7S/L3/42CO/3XQcl+hgTpo6rsCh0UEn158qui3PwKMJmzaCy1
wRYieL+6l6tPygZsD7iFoVVcRdgVXcmQZUNvBZvltydXvHLukW2Eklv5LL9JLDupjYB0osgCMlyJ
f8JNvMeJ7prCRmThpHXG0ImFX2sQhAAdAIE81ksIqz2XjAhWoTY8RMCOeFThy9XfoKGQ0Rwc+U8t
MQ7SwIxNp67PBBJo0bBcNHbmumSnPzo8p/Ui18+jtFW4jbZPTq1U3p3Iq7nvd9YYsswNppa4aE5q
BRBlPQyhVWPKBKWxi21czHewodYSoOeELjXF5K+65uVD/JPz/QQ0dg5Y+h6tVSNG2dYXQ8qHzUJT
e2p1oaahF+aBFIpBTp7ek6GAm5uQR8KkViBif8NSQgiiBEzu+ise11CdD7xB6Vh/6lNhK8gfd9qi
mq5hpvDWUjdkRrbVL6goXHKpMiZxiJ0WtSD2O/UnIMLjNHYRTRrcwA2TME1MvG9cwiLWiRj4Sigg
b06h+wCST//7XG6i1wxlhl8hiiQ8+z2g6K2Z1HI8NV9LgOlMtCHRBuimAZIsyJZ9/kJ1Z01AQtIE
6bivRyVgSCF38eG0EmzZdC54sWKzJWvQD/ZymBnYTwk8hMtm+77VJ6GJNm36MUXFv/uG3+h5/eTp
03CT5VlZiuR9SNaPIFeGQRwPBT+62Df1t0PKXzdyrWwuQi2KUE2hPabQGBFvFtW++A7w74M8losd
UqM53/uMb8qqYUvPJg6+bzl5VI1zjTDFGPX2EmPKExHDukNlpnjRZCGT3fFxtrUT2qtwjN0B8NyP
TKlTAqAVZA3hIrg+XXnE4uTipZCiPJOgH9hoFcTSRii/Da9J5iBhDjxEr5BxiVyjJx3n/tzPajwF
j3Xj0eTYnD2ahlJ/JjGN8rWAawRAJH8ySRR3N+gHU8N48XcEtWPYbXhngolUkO+VdN0NukFQC3C6
eNn+t/9BqME0iRRVTh1wRd/XwRD3ASjPDmBQVSZjkV5BZrxpQ6COKYAZque8y3HttQ9JQd3+neuV
gqsCQLUqVwzQ8lcuxMs3RUYZIBY0K5/0w0LwT9J+xXzdDoveuh9Nv6JM8iPfkqcLIYrifCre6Ywl
K8oVHOephwgRVfTrW9bYV8PeEWiXigXehOAV9UwqHkrS1LNFD/9y+xI+RgFwc6slPt8hCLxdXPKH
iihbin1WfZ0ZFy2OdHASZBXIY6xEdIdX5uQAEckG9w6PQR4EaWmfFp/RO0d0AgaN4QRCDHuYQmsD
d00RqWiChOSCDCjtQPGlYOWHT1fYNYmtSYCBDZIgk0nJzHmM4oAUE0vHzsZKRRLW+Pv1TseuCOcj
/3dxp26RFutm56mgGo3DFrAywbJT/Vo8+lrnYKbkPOurX8/ZQdGE84LW94rcpkBqMe/9KsPVcQZo
9o1GvZsTSDW4Fbk4tlZkJ4fVRtQYjMig9TDMi5ay7vIlaF6FiSl3UAdRZZ2cQ/Jwr3iXmwvx7MHh
1goE2BnWScDodi9PSUuDUGEMngS1RfjcaB1qSYcvVRNE2ALtLbDS1b0paxd1ElEUavand3/yw0c7
yv1USB+Q8hbIUiiuF3YogcNuXp99ktgUXL/DxRDp1lZkrDOq9vlsLahe3PiES16TgSSOAA6LSUJp
Sla0ICQcYUwtNJsJTChjpJv3Pg77K9J/75dLNXlxtqbraf80+TKCyvn3S/ANhElBDetxVU4kzSgE
joiz9+Md0+CYezYJLJohCFa2TSeA/th3lQQ1dJKkKzIqKi1dkHg+dOP6ArQNTdt7G5GuviaosoZh
o6ZpyAQSzPm2gY+6N5czZW9qfEQEyaDyiA2tGJ0Ee9PJbvsXYZ2/WKWnxF+y0fHTzLW7z5slyXop
ovyLd2RAH9xkdOpIrmCPWSl8RcrISZikjNXrLVgl0L8BUbHU0a/TU5TX6eZqQDLdc5trin9Hf7NR
mtHrzTs3qAnRsmOI6j4sf9kN2/4244qOhkU5pcpoV+bKhrzUVRjrNA0owu3UjG0HriuV8t0cDDt9
hUBSLS0ZsqAhKzpvJWZ7npu3X/7XwZgoIx2qhCC7+absVB7TpYGYWw0uDlqR4Wu35ptj3Vigplss
t7+krXevyTJm8sL3gqUNS5CfSwZ+YB14HSbODlr5aaBRRUsPz1hV6nLryRwAdtnDEM+YokQZtu/j
pUJQEgQXF24Sa5fBNsNCosHU5+B2fZs+thW0m0PfNWpfBOM1WOYNQc6EHeRYVgAonBZHwfk6ljL9
cJbOKkrnYh6DvI2OQb/dS5DaSlGZsYZvo8jUy6u3r4Ga0k/xwekMTIzb4LsunQN7ybJ8JBWCtVMY
XUzUGRY5wYnN9SP+sVmwY/aEO6KU73zp3p6NwvB+1tL871IJOFmFgwVEw1LUluTVSd2QFw/E8pEk
Sjdvf4B3XXSrcSgNiuqk2T9iFulRhKdIUids/wGtMeaYzxpNHRcAJ5Utvw/fDGxg/hKJd8KUHR+M
aSkp6tHLobwXSkhQ468qXUr+zcErQKFHf2zwDlCrrDF5iOE1r2ohk9iKmiieXznqmyTq229S4x2S
Uw98pE7RwAt1lRc/T/qGYJrA7bljXlqrqgScWbxQP//cg4ISb9V9F/7c/kbnSXbzXkVXQHXXiiuU
hhxsseAuOIis0N+CeQuTuwAt9m9upo4AdbNqlG8pnnvlDjNZcSEtmHjr4YrULuzaiRT5AU/4WdSm
sPT+FMFTHlEaUa4pqeU4pE0FtzybX49zKOKq12ZSeza9isddnQfuzznwsJEwvNlxf0mTcZ/utGA6
BQuR4BJYi88gpseO9W/rj0uiPXY2ASMNo7okx7MXLNvMkRIWVZPL3GLwDrHI/PBkPTI8amPXy3UG
HCxmX5JYLp/p5Hvj5blZ3m1kaRpD8jHFpXYQtFb5+tcgRBw4AMm5Wbydx2NfcnTyk9STQlZmh52i
ZUfYzIM0B5D9P/tLdQE5sw2Cq7lqCPydCP1o1V22LxJgqqWCLEp41Xz0ACXg9+mn4emPbgREHpa1
rd5BbKLZNuICTEI+sx5rfMbkWoHHPdIcH9cGWlo4GNo0c9SmLha65/VP39I1ireEYTifc60/iVS9
Busuzr7vmghEMuQyxBC9obg/uanpGnxEOte6TmGeUQ02vIUUCsgOOvEvDzoLpCJ3w/YsPw5NCh0a
nnz9ONdWIsSIBp6ThLNRJj4zJsFmUhV4qCoTvo9aRPkEqXkY8aZka6PRsoJFhtmOjzpEMkTOUVZ3
2TXAJPw57NHqZQshbyiP9O0gCl3xuJhVeWOE48ofb7wjGmSYunG/zGLSGv8oF1drynAqAEnrgI85
2Z9CKombPzs4gejM+8us6wHEsOc1OIoLNlg64c6h//KHvmKWdgYBu8hkq0MbeatYAVIgwTSLewjY
SogQXFWKjR8aagSSSc31yoTSPeoLSTIaXSJzEm3vwlLRBLnwY6Kq9LU4uiL/UPMhTHm5GeFGHiL8
XOgmuN7Q+1djfGnP4txglPa8rh7fcHRezZ/I3Bce0VSDSqtwk14pREoKr0CUxCpT6gzNf/aZ9ZLx
WzyUbNm2o2oKLdQaiXL+tx2pO4M2+WIaEJCTiaKK88WxT6P7nj7jJPTTm3rpGq1kR5WjDh/2dE5z
iqMnxnMkVCScgCUHILab8nbBjW1gaNtL9JC4lYtPuLY53q2eoqwvQbdvyr6gALIG7+PRsaVaX6Rf
gKORGTD3lS7zodzC80tkpicET+HF9hfBN8oKNYe5fiDDi+nf/vRKTE7wLiphYp7WyryZp5c04it+
yCzaSU9J6AJt8TfNYv5jbAeapFhf/XANxVMTkHXVpocbmp0yl5OgdpV3m2/FuEdlgkr1QxlvoptI
t+H/6AUC5NJzzpLkRfHzBptGEs6aWx+smFaNIaQAfma3b1+ua5nQiFeVId5dpHsP3fa2TbBv3b4g
McCXDuSSsJn1NmEBSjk/AcVLaA6EljmAmXZotdMABpNmw8D/LNVh16YvJ4oHIPS7MP59kqIvRUCV
KTSPkilN5dOhu/4StqqyycAARMI9g4xhEe8CCUJCUIKx539MEZXUcB1LObLFGJGguFT0KP4M0Wdo
r0i9T1vvi1yKv2eIFl9KG6yAJ1z/wxlwbE4CeFJLtWb8vQZDUpxjgEG01OA+o1+nuEWUInK3jtA5
HoHSZSikvZiXffNvUeYR0KdhnhY4KSDuFvyDIGN0eaLRWULsbbKeIi8cGSL1XhwwScTzSVOmanET
lkJHbkrwAZP723M6WbNhZCvSLBaGMfqNiSf7kZWEVk5mhFzj6GJZCBaEzpMKw2Q5fkrT96RB9Qgj
TKo67AxbjyiSpWTLm1UFe8O91vBlU+3nXUlW/HMI9d5n1rRl9sHrnDfSrnTaAzY7vL981XUBEeCK
nOIUsW97VfHC7DVoJokLHgMi8DXGOnQHuwBTQHfA59JcxIU6KrgHxC5eVgjfiHKdLftZp4N1mAWW
Z3RupJaZ1rYP9YXZduKbPObeWO2dMrpYJV7rF07D5Cf57Y56IItQdj6MHTlTflhvmpxPj1dlusFf
RsKGIGZH1FYFjWO2LuGux3iPfaAJ7s9oj+VmahB8hqvp8nTx0RIorqrsa3pjkEyV91myU859n/Bt
2lsIIohT8rVcxBS8reuzAHizNTi06uuYKENVnDs8klZXpH+KWeZW7kSFLqVi+qwuvTbCjEm543tC
AL4/ltqWlnLHK0ZT7RzkQCqU4I89GEjfUhIux/dmj9RsVY7hc1lOq7UyDXG6AvXfSYUzW8tHf7YG
WJoRRf/T89MajwFexUoA7k8xvyaPsJyGgHRK5Io9CeUrgosUhatFbl7oX/KgDMyfUDEU3bMiB8dJ
DZ/zZDxuZ3SvcnDaXM6hI3cbEhRsZVn92EUv+/oBM1I0fRQgZd3GU2e6saPaYQ+gImdfbaHNuwms
EbIbECk5tpk+M7Ay4UP3fKeDBbO0XwVFsJJry2jV3dW7EZ4Ut/nqi1jNuyGEeAQFEoCIQFVu8Pld
3hz63NSb9e+bwenMmPLRrIloW50j1NBCex/bIa5GXDv5/pZCzWi4FPrH6UVY2HcG+xTvK6TLZr1U
Nca+hfSjrspefd3TyaQ7A8Ci0PT5JTiisCnBM4nIXCHuCjonk7HaZWnqJ8OuJd3tRA8ObuIOm4LN
Zmp2ZP3XtrMxSxb+yDCtho2XXq7WD6lUYsMVIjfz7Gi3Y+LDwbCIbzPiZPdNQO6tlZX5lB3IR9BN
jV0zsfLv1HimIUWu90fgccKR24odsvZkhfy4OfJBgWOdnltNoC2uZzoc8ItALG9DU3eNY3HeR8Lt
DR9HiEYvOkZ2MWjKOCWsIBbZXUzgvJYST+mXx8FzohZUuRqxQHP/JeqPSheFC3YFj7MHLBY+BuZU
M3CLUSXfV+lS2Tb1YiXduGdIYf7ZpwcTrfEVeVey3zJ2JqK3dHliYr+3/vDdd3bSIf6BUKiKOsiK
jL1Kx/Bl4oqCSMGCzVJTFtgjMDFUMfLXR4cE1bPBeYjaUNmbRrEwN9ZuHWezXtBP+rvA2V3nhJGC
RHVnFGpvfbmuRUsLDeWn3mtIIPc4KAaCaVzCRNHLMfLPsw3LqTNxI+zOxOWuDNM/gA/wDopL+kKv
spdAaCxrHktYNesztLfw9wGWBKEBMrgd/L+bd0dlElPVcA5BnbsdHhcUHsE6V7r4y0Oetmd5ZEde
COBpQp/kNNBHiNtoTXMt/Vjsdepx1AAFEXY/YLFzOlVShb0HeFx51PGFW0ZM6ynxID9YBwY6g8lO
WPKFnZz0lJE6clxEHAS90PVSLkBF1hHtGenmjLD3EUACEPioIhuRMTA1ENWfnD9+QYbwswFJWzZB
kdOibnC/S8DS04tmm6HMgnwxG8liiAHD4qy+efSCw2C96NlM0Dm7GYybFsmsTPJ8vsiX2j3vxUKL
yV4ABymboFHZWA8mifhGqaDitKqpF6o13m+B7i9vU4TjIiPWHadrrRiMPFdVQ2AjMriVjQCyUf1n
wHntNGrbHSYZzvCROYaSbtAc4/1V1Polms1/4QWaBAHtd20CcnhsR3jnwgiR+LyRpYEZyzWwotf0
M4FeTu24Ka1P2oZV2G3103t+pH4briSG/OIlOc8XwufI2rjiKXXUIm8c+OgDphPnaLDiHWRVIBDv
nuoWtJ6V8FfhJcAwQXCPQOQAH8bd0EUydDm2KG88/hNEPKU6iOOuE7na82XjduDtA/CQRdM6cxiq
6hLk4QpwwwyY4LeAMKoiT4mMw8F7J0/sOGonMmoGw8MbDrJUeARjMC9XnD7ancnT4N2s3KX5K1bH
q6LNlUEFLYw5uZBNNGJ5XrWwSEH/UN2Z65fab6YxSFDiYWPs46LbbVDl8WnX+5NQWf1SoYIk++u5
RPLxc6WLIUXvBlT0+PR5A3pjzU+aNzUEunhOvR7LFCvkMvCcwvCxpFO3Cgn984gEIEnNsV6bKE0k
8flKq/uCT1Obr3nRoWFoDkpI+ovSlYaH38nW0Te9TafKiGhOKPFad1toW2q7d9paFGGHEIDceDYq
LtORAcAY91kdz5UO6xE1+JRJlkU6UohFAPgSQkpJ2XX5Lf8QUh7H2udOfBVS1dJ3CW+3TuEVzv1L
NidsYWBuwqW9+ycxoTXn2sOsLladyDjAHWVS75QstrgL8G3V0YtRCPIXEBLu1QTmT7UiAkdxnNSu
PVYNUm74/8aH0zkQz0UX5jLTfLvPXZVkHxoOmpvtBuD+cMEZItVH2oLnAinUWuKEsnD2SMfIxoxd
LY30QQFMok3KskMZvTaPQ2mexB45WIoSKxhAhumeNXovOoBcYqVg4r/Wet6SbpjnCBRy0ijqM15b
EdtrLTWEM0bX+yVrQgY1oO3+7sln3SheBklPU6Tx1tg24nT1HFOIy87MUK1xkTYAE5dEX2H9tmee
Xsi4ncONk6xbnVXRyz8R7/JiBvJN+pEwCBbdJ1xYFhehLhhWcoQnTGdODZLzmwLeiSav3xDVuFfW
arE16p8KK+dCjXkiyQjn9gmotGQtB4OVY+A8JPw8w3M2MVClRzApHBkCmEixsAB5tX6mYpf++RKy
9U4aZlceNv5fUFzbdKJ+z6aHNeLYbzNPk/WSyqJagSfJ6J3A+hfB0qX6+auHWcXkfTvX4yoZwz1i
GGd65Isj6vj2uHiTBv7iEd8N0rzobZ4UlDnN0cMeTNngvxIsiDdPr9Bs7s708lR6eJNl3UE27IY2
tPsK6uB9VL/6kv30V+fc1+WR4tLUK416gkMH42xD5MzNGByvALyqF7cYxsBfz0UifdRU+cD0FXCH
rLUj8qxetRjiGKSZ0JL7GChOPhJT3zkb4c0q1VAlBsyxSk7Hrks7/sOFKxg2UYC+0bDf+3XNkN2O
gQaTF4Ho/eV7ObStpV6p/pGnMxveS/P/1ZGb9ZO3zL6TvsvY3YTWUYzdhi/Nf4VOJYseOSE179h1
/a1MnkGTFhjQyvIbbrRh/Z2K5pYtXL9gsMgP1388vC/VqUrj7qyLmre7c7ShLsoQ8bAs8cclK2za
Z6BSZeu3EA1DtQZifOIC6G8qF3+87UWMh6sBdI1LSkLH9MqhCtI8VyozOFcWIan0ds3zcvE1xLq6
24ZBLJhgeZTW/fS4OwHTnGRKhbVRaXcKiOv6tnj+7ujso4DkqtZY6lBOh6Elu5Vd5YOy6Uk/0q31
mYllKoUhVA8MQLsMIZ93NaEND6A4o05fmsOwsV9noku5/5xp0rPR9JIIopUqN1kMPO7qE/eMcH8A
wzz05w/t6SWWL3pMWy81Abd/MjoaELyTQPFeT81ucK3xNrPtHuB1p3T5QXaXiWEUK7mo27BWc6BM
fLiKD2H0R8Twx6nEj6AFIS4KejQ8PBfVtXbUpCrd3/GzWdxHXTvl5PRRjy+RiwMWKsVQLx1EC87v
d2GCV4sL+eJXsjP9CDj/Z/3Itt92357TaOztqW0m5XkpPn4W01inmd5ZZqyW9H0wlT9FfnSSXeNC
0iJAGqhfLqUdsUAvwjHwnanfEsuBKsaaddyOp52i9aY9k2YOr8kmkXPqZc8R3mZOmyvA5JXy1f6h
qywvmf/6tJDgDXB1oLoHwCAxZvFu8gYxOmiC4I+BPpFEmXtpWAfWpfTAdqdLBzI2wo6BapVNFJLX
VLPeqmIg/Qlg6K1k7SG2ZwTPUgifQQKPYKBubD+jCakYx0aKVIinbqB3U5ruKcXs19oH0yn7us06
8sWYDemmG0AlQSnJQBz3LoQLq4J6S0jxEd/pRF5deVV5t0KcSI1wJDaFm+7ZlpPcxBIKfp2CfA9a
2rbbumHkSrFoiUMC3k55CUHYHAhrSCcRzkA4HWlagWP/SWdjNeO9qfXTrgJBcH/qG3pELojvniHP
YkQAbCxHn89SQ3bOWAurxClC9M5iJfWypgOEm15M8kVpPLbAsWg9FpLIV9q0CnVwp12m+Z148war
f9V9bMsXHhqo6rTMuZhEEEpoXNuuiEtcdKhR4HNwpQWEZQgb9wRa42A1KefC+PQFOOgXzr3ywgX6
jeJWrX5FG25Yf3N8YzyFnhumWkUQe+TqcA0LNJxNF19RuJrjEbNC9rwWvgnka7mm0UFA7gmWEo53
N2o7rgoPSYorUdhLcNzigMq8ppdXgsmhDs4h+UVOnsGyHWpZ/yoIv1ufEhBKKOK52QUGh5YaFV4J
3PxQMgQfBai2AsP5drDHTyRvJ60hiuKgEnZlfYHFBN/N8E+K34xE+cq4cVHlafeb6JmILzZ0DqWn
lW8RbK5Z5wiXDgsCFOmI74nP5MlOI1KgHdsiT9ThL79lYuVuApoBxxXqJQ8/TEZkzdySX7kkRTrX
btDHafDnnP4ZpzPqs+EQoAEXtC+Wwqb3PVMBFCNug/D8QLx96YH1dsuKX6j37jpWuIZpSqKe6gXM
y31mDF6zxR7HrEYVsOqBTstrtnNFbZvhmZoBJGWSkeVhmeGW0d55phb/qe8VAE509Wr6uICxj/AF
ZWQFH27mMrgvugWyhRRUFNE4FTAMpM2UY7zs0ARPDE2SDZ+MiCNbocTngoPFD0/Ve4G9iIBvGf89
c7Bl5bZUJaNcZuPrcNnsr75RnrrQ2cnQnsyrq8ZIawZhWUztJ4LUTy3xqDFc5GuFZUFGqj1AYCBz
jqbesmJd9XdeZUdhV5gfPojCJzfJoa1Ju/w1kIWy8qeDgjHk+SoWJarKbwQ+7HwJ2Ii0eRvJoh5k
2auXlHif1Rmbc1jZ5rTNW8yU9WN8Fh14eZHZXeNYPLBQ448FudgNAPHnWWf0m0Hupor2nSiH0nwg
sU1J+8cLZcZ5vdWPyrmw8ESGsGSZ0D1p0hHFEyxy8mwNeUqswC03UfUVKgMKox67SL0XZpiruCHY
LB2rkL1+zpUYoot3R0WcvihMkLLsgUuccTaoyoQUxecHmOhMPNsMcr02pQDqcQ4Twf+FH8O2XrUk
mOhe1qMPDRGKzTDc5QehoVV5BBpZNYgQcY0Ca+ttFZixBpWMt7mWrJuPHxedswbwUZBUuwSlnTZ0
7CoxwlZFgTF8ErkQRngz4T6vVAJcdueiGnygfVgTPa14ZkmKjbw7ke2r1Tc/UNM/wavgKl7r5bpF
rgJ6jbjeLd/hf4EQYv3GJNxk0WyuAP9fbXT+SJVFJgIjv9AIQWAWaSvKv97otj/+Eb5Qse9sI/1j
uaDWKQ9A6IRM7b9dbWKhv5fUdoHRJvc0rl2HzUX4Nt/LTfYH4txwv20nratx8muMw2HEshkKR8Jj
iyobOtRe6MCf+TudVG8u5j7ZrO3vc8bFFJdiusbCgHfuwwnQ4G7z2gibqLWU69kQHa2zKj6+Clp8
DIjg46222YRP5NuBkRhzhA8abYyCFb5UZYMXObIvC8o9kQ2XJeOGlpufpW4/UDYC+j3qGhcI9s1b
CH2vLaLVIW1IQAHU949enGiLOPPTvIqubFH+Lvp6z+C0VZYivhcC7yyB9qW/GRxCh1BePu/A/w1K
QdypkofHURbBCowQ1mc26mmFmszlwi2LYEuN3YE07A4p+g4Y+aypOVpcVGlbiaZx0p9tMeB5+uCh
37o1Zye/wuXrEbfUToqoZGTim0D0GnNQQlYC0JlfBKPWFSea8zu/abZ+PgB2zfK/7sWXFg6/auHG
cNxH7iS01xEkguhBIJpOM8tYzkZyof6NExPtbpiB0TJpl+CRDpqt2+2Zk7GcMAI0hbBZrPclCdnp
mFEZrdkaKyanRe8w/tuExzBc3Lk8wSdz7yHkPul8quZtBIejdY32zYecilBb9OOzYq+GWuwrrg0g
3AlUVwAizGosu0rFWO+gnPc70MvY71vt2c46NoOJDqmQEsIIQ2PWBcitXtW/toRaWqovjOMUiXb+
H78GjioZuLH90eLlWm37kpuxbsFwdAYQZYHC9sHKtKp7EI9R8MR/HXS+D6FcejD1MOWjIkA1x935
nfBnbFB50CpPrlchIuVonhS1HRd28FhPDUNUAcrc/ZsQYEGpVzAie+v6zoyDPzzodF9ysFml7aTY
VKfo980+1oCn7gjQqGV9fEhXDP9gMv3KXODVHvv5LgaI1fWRooGYNWcjlg6tXEFUsZKNqhNnsoFB
7WxJ6lmUq9P8bs2XiH2jfUwLMviAnXWQYXUEYMHzB73hI8cu3OhNxgnv0Kua9ZIvEDDrHwp2jXal
4zj8zlYRhZJOajhJDQu3Ohlzu0ns4LydflcPsGz2YIuLy342/VAydD79Y9nXlRPLw7jO7WuJ79jF
evOgFdnmKfWaSfGWBeS7QFNcEIhtHlekxNGXyC0yKMKXKDTPrO5Ady4G0ZqiqrD9YD6lrSGqci8A
4JtNfrOKQg7TqLRNSLFyzNyu798zQNgBkPhEim1Se4OGmZs4UqXqZZh51bhUvx7OY7Y2H1tB0P4A
ryRPc6Nyw8Orz99pusXsNsR82IezzmCyuuysDAyfUpVFVn1iL4q99JwdrgaJRfAqouDHpOai9Xc3
civLeIXIMzt1ksgYy29vc+vq1bz80zacXCN0xMTb1xzgZqsVaE+/mnpHLXsnsGmSBN62qmyeFWEY
ic+66/iDj8EtpalyPH8pyzBsYRKcMDcf+bXy2TspHH6bJI4u/+Ytb6DsJVPSkkVPheeePGtxGcxn
qHi4FzF5RBqD3K+OKwZruBn4+qO6H0Uaz+ECoJZjr3uYVJ3gzpnPMIJ6Y4plpFdycd54pS0dNzRF
c6HGxfSTvvlwupY/Lfg3ObPNn7e4BtU8pIR5ymJHTYnbET0jlVYhL1ejbMIHcFXoC0wwoxWashL0
siQiPU9b6guXaoGddFtbWF6FBH0hTUy2lglR8MdBRVO1WuPS+IDRdKREI2HCak4CTzBlogxsKoBE
S4zf7m5HrBuncbhpHGtL1Rz6uwIRnciqK8o0dhXaZe8s5IkdV8Oi34x5x6IhNbdnrBGFmCmFJa/H
EzRjknzc1lzf71iaCxPQdw/JYaeNfLVX3RIFnl7MGCXNu1ZMq6H9Cu5URx9+8yLU8xeAqJZ6avKR
9onAVg4tkntFkDA0Twq0Lc2r92idfkKiZ1zH+9RHbNYGquknzsncnia3gccCF4Num9/3XauAgyme
wc6I6N34rCORa/OC9YSU0VYwvBLOBPSgSUfOU+mUwxpRXFbxoeje4yoJOEUpayjwJWHxHTQvL1LB
l5pXlrzBc8YGVOojTxm/x+vhPf9KfpLsndkCDNG6rKh8N6GO6YDNhNky/5MRQRoltqWxAk7iJ8pC
fBibDL46UmzNyLOv7B6R3e5y92qF203dHKBg2AfWAU7k49mHTt9tc8OcUnyO5pBCaZo3vzG4RCge
oSEUo+kbBbbsGi66jz14pRMhD+szLtAleiDkDEzZss5crO/1ae0PqsX4C661nwPWfTUo3j3zLinI
F2PSLiK6tcdzFvIJm4784IeukgXyB0PMTuOexU5Y79eHsyUlgznt+I0cI4j6C1cOBUSLTJLc0FZl
0x5MO3AnsMEYxsO7zmpDSLY/aSj7LFFU0YL4SZJNhQEqfRfMzP5SnwFnhx/85uHWoL6HfFo0Qst+
1nPK6/0PTIVjZBmHKoe7wSrM/pUQquzqNRUSycTyiwo44OrDryBEQ2j5efuGq9eshdLX1e72x0tM
CLJ5vwQd7x+C0teQt1F2q5x3UKIeZH2Z0UWHzxENQVC2MecwgSacbDBZI5uYvAC7+I4TpvE2a5sM
hNe147fNGWIs7gCSE0+pq4L1ryCL69Z1NBxrtk8taTQUTqkNA7n063Lgr+yUiiZ+jghe3K16CbZv
o4iI5/54oe7B0FecRhf0AxKm1MaH/9cEh2zz18+t2pGglG2heRpXxcHTOVSUKP33z3kXmqV2rCN5
lNW+DbXEauap2GhjDTr41tyLuCNPFaN5Bhd78oKMkwh6TfjDOwHlFa1gowe7rVt0+hqa91/vH2ee
BxDiVdR80ydp6+Hu9J01jo17TFsgPdc+EC/KSA24Kl1ACbSOv29BQI7vKtgC42SHCjr5EzgITMYx
5wcqZfxAX1I7Z5HpkV3o+QEQ0nE4mloriagLxtb5QeHaV7lnxgqpacCY+SInRNB96tuD85oSyaKx
+IWY2PDjuYS5WTL/JqprLyXXNJixl+VRgEa62XtWDYRNv9Hve2clsenffEVIsBh52Viz/kz3nmN2
X+O1T/SLh7ZOYVnTe/XgUFmLmihmd2jHCbVhlWa1JjGqgXUESHEZBqdJPOd5ymIjGhuBBNpW9A9i
vONbn06C49NshCVtNsUqrxXu1oPiW1HdT7TxFWz/G6bfroCK8L/+aVSKNIdgzzpoGGU6NqvyLSk4
EA4gD7ptdYuL56w+eKinpdAOQJAviKn4qQAUMnGPtN8hLaPu9YAdS/cY7mkDvuTXXXfCzLJ2PaQm
WPdfV4L8Ew6u+/6rhoIssu0THaiLGMmG8A27kHV5Sxf12FKq+3cfUs46D+xzKsUB/PtYgoUCuM30
WXcIc8kvU3JPaq0OZH1ujonyThHQrKZ/IP0b+suiNfTOpgJxWJsi8kCO8vBuUT/x9+w6ZwOcf6cc
FzhLv4eM5Q6naMjJerC+2XcY0awPLE7ypJHF1UtM2sn3TibG9xOrNPfzgxFiz3T8JvAKbcSGF8Uv
A3i5b7Svx/0CJ1wP5AgFKzhP3yijqpy8YF2WBjLT20xRj8HEPfH0782g/i6da9wPyHQoV3XfnG6v
kAopL7eL7Alj1RLX1NYOp6rPsMejLmskTcD+cPtamOnYnsJ65cKG1nDfXCUTxvcf1lcGIcw/g3gk
jfjhdy+oEUby4/947EIob1jLkmbIUYMy1JkIp5gyISDGCdN54dtedNEHV7vopWo3LymbLO7gXIoO
PTuTC4eswe+6lpp1r5rY+EvhZXnB4/uM1O3VSmvMOSP0u2UiePFSlQlGsz1WQweUKb0w7IWsfgcm
/RngMFASorHDR+05HZQNGBJlWzNzjM+qmZjouqypTw9Aw6hTVSosCnj+epmbsG1Gy678/SvSOid+
3x3zmFElFQFN3/htnfAQPSO/BV4zbZwop7o5y2ZQVhKkHAKfMIfwICCgGpGt7kRFJipcn1jBUTjR
TKXSuRg8tKoTnDMqKuNz0oAyaGJiy4nizBzhb6QK9wRl5BQJBITf8GLg3IuBp2Hk0ZcEUB+x3auW
SgJLWjpbyfXjgpGPAl2rgMLxyhX3+lb9UDeYNSXih0Unjic5WvoPHLbO9cQI0t1Yx9Agh5CBURxo
ZOLt32ynsyxSiyFiPYpPx4kZHT9bXnsOkPhH8wRuF44aPsKUiX9vi445qw90+wpXdGCrAuz5jxbW
5orBdlXYYU6Ek7D4/z0utKNiwHvnAsW7LFprylK05Bpjf4q+TO6qZ32uCxZqQKgdf6fGfdcdQzEv
D3/BdQ77avyuNohHwIN68pMZTPSga5/M914G8r1V44TQksb8S7qj6zZhfG7ryoX6QnA21ixTByRM
f9m1RRJTIKLuUrJ3LNsbKFQl3BpTHiIeQpkiC/kEmKuU5zjcG2Yxv3b/jg+T3mLZJ19alsU1yHum
RCdvfqZXKuxAnYrej9w4boFtRSiXTK66k/3uQpiiQMU5y+wmiRfkSpQxN7hUfRSbr96JfFwyu52g
4+qUEVZZnivS0x7f7Jy0k3SAbrsq0PnlxtPrgUjXWXjP569tpQIZv7UPMkglaWOqECGSvRNQvfmb
MDPb023HDkfxjQdczJfSy3fZJM2bImwK8p5yfHPUHyfvioVktejGuggaF0BUJlEfsbRHq4jc8Rzi
b98VdEjLnbl/WMiATahtDrZLN3+O42zTG91XWEmkhQTX8MnJoWcnDV3J46njKW4CNpOP8ZZRdaw3
qetQYidGi31sUmkHXBhOhRAFnZbxvZ3yNNY4W6VpkgZiyIckowotFIzl1Wu27cyG+q48/qV4Ybm9
Zl6mIq4QvtL/2zI4j5+OXVumeJmYRAczGy6TQs4moOJcaZaGoSaSDK6UWXa8pFgSB6QwcjO1S0Gy
0ScEMwWoOFtulGPye3ylDpt8Sf4bY6z6Ki7OujFEeni2yFzfd83UKWH80mgT8sNLW2PoohPhYD1G
y+WSYwFF06xBI39nkNEYrBWcdSth+uCREg7+HxpV6YpekxWK111b32Gzw+OJKHiZs9B8ErEofa0P
JKXasEIVXmF1KzBsf5gKyoNmwAhD1c6fBhsvJ2PFW7cyUULYHARl0whe3kx/1wzM1gNM/H71OZjD
KMQbBgMS22H6mFR2aqCo54rCxxzwCqhN+4mbG43gPMixuQyv6dPnZGl7ua/Ba00Thvd8E//5Ww7n
zyfqudY1JV6vea/e1CNoJrMGpsREyDfuRe3RfF3cpAlAVsaGYfjiPzZk9pS5wmMOyrRRE+AfzJZ3
0yFxaS/WBqM2G6ICDrjGMwUbRK8mQaxHa5JKhZg2+t0K83y1EXL8cLXlJtb6mp49rCNAXWvDNy7T
S0dnfce6QMNYqj4hjlQfDatLTTnnd1Lo3OlhteDKDnGlnyaI/5jQUIzpndypba/gmLk+hqMTwGGk
fl1HiOb5jjY9oOPHluywNycRRu4DaC7BDoeXocZ+6MjepK5jLshNVOcp/5JdZe1xK93zuH2Ucqrd
yppeOhNa34Qv6KAbAxywbuuM9dERfqQ/E2ULirOZbi7rZ0mgZ6ocupf23pBkyZTMdNi7j8eCBbSF
5fQk5OWNfo28ycxEcJKjyGG+BUEt7u4DHRP8J6cyxwT4ZjbuOOYNKqENruPYiTpVyGaFkeYsdOOH
UfCYqMpMgPl4251t1lVmXK3ppQhtHzqIrJTfgwohZzsf8AsrkV9mhXrQ+YObSny3WqJyUuLQeZ5f
pteC+pWsxodl2ggOJDiurBlCYICrhWPX6y5SXzuBvNKnZ2vlKjPmSamzue1cpR5L6sD6DJWKewaN
A1o1R9uDsApK6cUd4i9aujfK6E8cE8UORjq8R1L7b/ajHvlRyXMy984K5E+FhPGTXwI5vugSv9hb
Sme5+kUe56e+l29lciaLbFflhlTTN/puRQcaSMd9jgld0CJkdyW0PixG+NYNuycw55LlDyl1F59Y
EwGX6DoVOLnC/hyuc2HuDw2FEgT6RLg4oYBaA30pFqGyQpAYSMCYVH8tLIYoCZDKsAeAQBtMQGhk
T8NGK0LzfG9Vz8Ecure7C9tnSqy1j7RhK+3gBqHnxQ7y5flSV5MSLx14XH4zhHw8eoaWKG5IguQk
D7DcI09gjPmRzARzJv2ypOZXd1ykHohHBUxhKK7Or5+OEo0Ngesx1asfXLECL87TicjDQu1Cbtg8
0WTNPNWcjAaQSI13bunUrztOP5Iu8S0Xad3d86bGL3iOQntV8LitNSRYHtF/k8EsSWHvTXIyglTY
We7Xl376M/tJ2ddW+A5byD1gv1+aqxPcH0iyqQmgHEHkk+1avrOWFK+BKBmNky6AYiKxfRUbX5nY
ns5SnwDi9cl+RGybFq3KFPs42vabEa2LwRbdBuyQGMVkuKnhurMCaO+Sjc9RkalFIUsu44dcpSxE
65dKpQPPzOeFD3lw/Z3JtJ2JiOwyQGeMnZUL4mEDZ8foaLMJ6NqWqBdvdDMZAkP/M1mgSUTBPsKv
KKLSqsWl7rCRZkD9C2N9yHhp9A9HygbSrW4JcoS+540S54L5e+aCsGKfM9NdxsO8Dq31NeAONtzt
JbVtsiBnRUwZpb9o7m3R1fPPwSfgR0hLYQ0znX6pyOWJOLL1sl6Fe5V9vGJVx0oUDFbT7gcrwziL
w//Xmn/tIKB+IsIQfCV96feHyw5u0EphRA7KoZDXni8NILVHaToUaNv7kvwf+PbBIPxLEevpa7P/
dpd/yv/HzDtetodUFodKp9dwxvDaqNOXh3jS7Fj/3aR8YPyBdb/hU1fO76RvOp0ZoEcwcugA33Qq
7Ai4vlgOavjk4AJpxd7YyhiyGixsA18QTAdP8LTY0TUa82LvAb6g3vwJzf93uWqrrtCuI5YHf80U
BBX2DLkcIbWbY1Eff8VSKSlmg1Ut/tEh1DclEW4sXExS5BNUmFgKSPPw3oSTeKpKztfZa7jz69t4
RvzJOHvGOP0RsAr7nZcaNH3xBxhAyfRWLTlQ3mILs0E2Hg5n+PckJRh/PTCEExgEK3xtzY8s/yyx
RCcG6uJSiPfB0ffRS+Lv+Y6m2UVQ+6Nb2D4mxHLhAsBJ/jMlOc8rOABebW9AVoIrmvoQ8Wy8Lb4j
MPsoZ1pg3gRayJ5uJCIz3YvtDcUNSc/vd1EGeZ3yN/PCb9Uj38DZ9SSVtQZIC3qppDlxxaZb1Xpx
OSv6BVSq71Z1041H9IxaPfXvraMJdyj+//rufJQsMlrspNeJiMYn1rddYdF8XnxASTwtwfuPHo8B
MKJdrON11TJZnCGdRSAU1cXGN8pNsXeaR5NXpKdhgVhU+etCYsspD0sOR+OHjOs60TJIDtkU9UlF
NcyfvIUzMVa9ETUSpw3PUCHN4jcUtuhRMKi+xuWh7nF04IQYS3HFYEyLO0YxrgkYyeY7pxqUM6dE
AMfn/VRDAdo48ap3HnxX8hjBnRV9NQg9kwkM+IzADky19U3x4j/phPYUUY/J0wYgAAOSvKWnL20K
o67iVP8K8fwB7/Uxxp/vAnegOjHGkD998Q65mnPJ+MTGpvzbASPwtLRaAQrxfxMhomgtl4Ta7pUs
ppbrZtKBIfbtJF5uf6ikKhsXMbK8AgR4lZBa5HZOjFK+3LsZkbbPmwlL1q/pZcDfN2C3omQOU8bH
3RM8+okTTqtZFJtSU9f5gCh0JOWuypLZq3Fq6igVGoXRmZAaB7hHvFvVwo/AclvGeTAALBfnamoI
aXPquSFhJxUdjGQBN2/d92sG/KJGCXueXjt0nkIfEa++Lei8TSV2EmWen3AO98fRFwAr8V8Qvibi
faqzRrJpnyqepFOCBvqK1gQqoyzUhFcSw6v347aTE2SMpv+UT2tlO9h7oflPEDU4Hm9YDYadcHAI
wkHATgu1tJ4Ki+3Tw4n/g1JZ2IiayissEkXHg4yentbVknZhIMn1nYg9si4Hy6zlklzOZWRxD05D
lMgCXLgcY26B0cOcvp8F7dmqnTxSQ9hBhN1dB+OjhSNAvT4aJMOpjtfgGWKlpXbe1mBUHVKCM6zR
qOVnVBJnI56cMJnIYsovo2lrf2EEyVadH0suu+oQTe/dzfrCnqGNJBdXDjDx7KkY0LukAH2csHU1
mRQlvjqJOMK1dpZYGbRcWO9X3UmmwV66wj7YSbbTl53TqPEJvIWQVYByOOew5nems5f/TN0Vb6zO
Sv2OkzODjfFhGRAcxiUKKl3QFra4QZfdx+NxsoCJZXYYK8LQeGUm//DPNfOffnGoNkLnhgG2gCDE
mKvb09E3C+HtquUrERcDA+JqR/5RRCllOSKOJYXm6Ahmdl7BJIGmkWaBCapMTH+GIzpdF8Zz2Jzd
/g5i7st2p0UytmENwLvKj9xjHSB/jUcvULwYKEnvhudv/2dmsb0Avcaj9XtlRHNEamqCgp76FcYw
hmEOE82DfP7m5X8L3ssySeVJ1BidvIE4e61rTwEOnvjSIa2xmtSAlLxZsfDw11INyxUisg/qFeNW
qDMKW71GErgKX+Kq7bRZfPRqaGoihV3G1SQpb6SMY08AYeYAcGvGWTnEyCImn6eNp9LOnPs7XoY4
+b2z4Bedhf6c/jTZgoIsVkP6Y28eRNkos1woPIb+YxofCX7yuY0bGJK6Gqt4WJEB+6+ps/aZv2CG
nh7bFdrIBV3mDJDeRpZd+Gcvat1Xr76kSPsC8mJ/C4Yj6oSskK2I98+iLB1QeB5AxaDBMm1FjcJQ
xXzenK0B645bOgQxTM6gHOfHRgfG6TM5zYqN/kSwD2Ps3UnqPUgJO5Lsf5vVpZ2W0WBdmGoyj3uO
45Bx1OrLHLxy5KIiYb5/v1/K9Oeii43PIX+zbHebBoyA3hyTHUjHaCIDcNRsTbXOyWAhjHRtFmPg
M3f5/W/I+extMr5+zf0L8hjznuwyVKLvaRsQsysvzupQNAQKwhhaixLVc67882PQNvXHZGCn7+L3
0Wz9Zs99W7F00HeDXiQ93EwCJnx+XTc+0jzuMKm1RdnJsEIBVaOQX4uxCnd3hLf6Vg9RkH/w8QgX
Ol7pi95h2GmyBQpFhH/fwtboU0HrPoQ1PFNqwA6WVdvqh2yORIA86R3H3dghw2Q2g8pw1PoNtEdF
ZCj+XEVSY6WOUYU31iFXS6zoWtqioavLZOoOnCv9nw1KoMaMdqTUUgMu+BZuJ9gJHzOEpVYnltNj
yZ/GLoCTa7ltbpo4An8A0AzjjFiAROKmwKBJK0Bg0fwYCeOckJUMDkJFlOjDiCQaq5gMtaEYqr4w
U6MgmByZ1WXxGaj3UVXt6No2sU/+/2KK/T/VLzWsso+/J6u66gXOA+tj7b+xd7hhaxP7/zIs7jI5
u7ms9dGMo02UD+K9+lnoYOaujuBw6IjlU5K249q+mF8GqWaGs1/3eg5kFQZSJLmE4S+2AYmF9+bW
YbhW8/UroncMvpVcp2LPwWKcIHJcu4tDe5yBlL6xFCcdZl/ofYvdwy6EK4tusllQXmoJNxNKywOi
VnzJrcFnTldyHedxWdhJK0+dMePYlfEDGrA3lOmwfeWBYXHa1J8T04I1fscvKn8cwz1gDsgtbpii
HUmFkoojR4Sf8KaGnfLnksCBdJLLt6q8l3ygPED4fBST/YUEQ65ZDtxsAue9gvIn/SGhNvqxcsY/
2g/q+k8doZJBhFUHWajhOSURAWsoB1UgIScJc28Xmhz9W/6idNbr7QXgYlDxChQI/VDoVD8b3uLY
Isp4P/4yjLmzhVrY1SFiS2Ic+62O1pFEpCzxMjbxeTiwM8A28/kpiTNguNxUJdoW1dH77629XadT
/GbZ4XTpS3AZjFP3kMPiTpSY+BTz74q7de9rJRH6BrHe6M5Eu6yrHcV5OiEolvhbY40i9KIJjsES
EjeXFMCOdtQlSwVcQ0FiU32nxOSxNReH8sBR1k2U5Qm2Rf3WWOMtccqU3pZjnZ0HY4k5DW/w9xhE
wEoWJ6//vl9UVo5fBoVjVFjmSo+9cdGYI6FeMVSnFA93sY7QzwqfVnI3aCNp1D29GJXNP91d+7IH
JzmZ8551Ifckz/GM20EXWzFUPOyLAzR1iEZfI+4w/ze+t0eZrZvxkOR7eAP7auhqhxDH7dw0aVbs
UNdTxXu41k4P+d7wtPKML3lqpbmwtGocGuHEImSfDRFKkCTAGNEmsB6KhRn8w3XRyaFS3gLqVBs0
wRzRRNs+eAlQOFeHQ/b+rg72ccGx38u2+ySSAlmUquogd5V8CAB5cIfZFOypfHz9CylBu+YCUVrP
gsNtGAKbnclKlfOKlef0vEU+d2yL9YO/QYtWcoVE+qQSNHKwiR90UVLnWcqVOWF6p0aroLyakccX
LOyLPVX0CIWlXa5r48eONfa8z4O1J5bSCfiqyXAPiN0JrQhelWyQAO05pSIy0MugMWtLmLtrqb9A
YZ2D0Nfe0bvFGIP7RlwbRrWM7XnRTO5G6XtdyklpUPafTQyK8pUbdSxhJTNv2Hj3aZVtBB5bkpLV
LuSYn0L8PEdH0RABYeHnG/lcg++619ASUsH9zyr7YTkR0SvoYt2N+zyrTcGBPOsCd0WPS17VOaTG
uwSCGxFmxp54edkhah8iSL2gmraOxt1jhGITxRCfNx+t5cPEGOVPuJvF2yZi8oSyES4tkbNKFcF8
s26ASI85c6ydkJGs3S1o4ycl9lkUgblvv3KWCBvSNMVaSCfvB3R15Q24jL/P9QlxE895hrPwxGtD
iO7okGSCKRXTmKR5yUEi3gdG+Tg8aWtJROX/jheW1kUOc77I4ghZfEMVfBJgzpjLZNT2eQr8ajg+
5cV5ehNvwNQmr6XXqFixa/mmYRDpLKvvgxFPSSnw+ciZw84hUlZDnbFyPRo1sQF+BSBt6JBb0hfi
w36LR1wcgp5JtrY1c0hXZNKjrKNGMijria/20m+1pUDiW8qM42AmC6DyM+fJscOvQxfVvWB82zhD
jiDFMZsngGNXkopcbRN4yJfZVUSrM/2LzH5gQOYFVDAhhdNmMUfbKHlyqERPsrdr5QOWva+W0tBr
fHnDaDPJCDdlRVNDRTcJSZVY3X52fAG4WYQh1nbDlRE41+Ax/M3diqIqwSGu/H5mev+XqTxA+4Bn
P2DS9IDzgWyxL4YGJzrnZiF8e/V1RWAdJ5q2MN2LjG7LfXnAiTc69PvcMqg3msQpQf+cKPJioWwA
GKxmXpU2Fk9dQUM9MssRgQTG0p9xevWxJzHR6BLVIHq2o6Zg4Ul3uVN9JngbBIsPrRl31fAkzLmi
mxOKBWf5CL4ncaG/GNdidjqAIFP8eJ+RuXEniVVmtwVp4UcekbV2Ikt/yZB4LukHwDTSjSOBnsvj
xrFQm0Rnzoy1uLHr6PTb+qW5mjKC6N2Yad++FxTxoWEHm4+TmGZMHMVsBay6+7jwxvfOQOKxLVFB
k/viOnzPZOu812aLlXG+AlRLnxRINWB1KLijMZRtTKgvnohlVdOVrdrZngdDGeSdfLTrqeq+sHpC
QMjLquPXxa07hDeAG8WAOqgBdxRa/LOF+dIuOQivXnkjjuWnP6e5pXGCGHnOLLD2zgalPqpZtCD0
SQUT9R1MIFCkDD/TlzWQWmCoWewmyb98+OfwZCakxbX6UdXXAxPcH9D7gLR6y/ud7f/nSvaM1DvS
sw+LdZK22TBAPqVh2v0Vm6Vom9HTjCPnNlWOSDe8c1X/B6BVttmR9sft3OfLC9FfCxn1MXhuAV2I
tVsYEuJnkva5SHuxHnnBOdzZAPWIES3BkNx5UvtPVGFrL6Q4Z+B0MWd/ANFnZIc22GnAq+hDfpoc
OzAXvsWuf4FFQ8coCzlpPPP4vJ0BS2Qi0Z8L4yFX1cZ0/p8ZvJzuwpP/kMkY5XyZFreqEqMMwlh9
S8nB4gb5pDqxC78gmRivqxWR4F+24gyFqLW+t0JyHsQk8ymXL6Dl4j2e3lFCPvHNz6jqhV6T5XHg
G1cvUkFPG4nvJvc+pqY2riVrVDPU1u5QixXhlMQgWs/f2T7W9y258THtsj9fYg2I4PG4cqGyVuqz
+JihdGoqQsoopG9A5V8lb3zWyIiySsxZtEEZCwkORWzEu9oHTgFIBgD6xUHWS3ol7JHxhXha9ixG
SGYhoiK1A5NHrcr96U/9LJmYzpgJeuOEEsxvd8dEhVJm1ZRnsiJT+5OaFjmJCFsxBxGAFRnU6w25
+yrHJROjE3OaarOCtKL+0vDYU2KuqWVr3NpUgGpekNZuufjxXyzwli5cyvWuOQkdd4P6GTQ7YszZ
XykmGj/F2czC3zeZv0Bfzt+JqDaAfEpwjAy2hRpB4fdMPSKLTz0NlOloHhM4vsx4jGfXDTqt4vPW
ANo2KUj5b3jgh/avYJ89GTcwIX8SXJUS+WOPu91z3H2EryzunQP1UP5b2PKlRi25FdhtI0g5Q0OR
/8CYZFS0t14fVARhI2XqKmTRTD9ToiJYHfvVzZIVBd2I36BSkOgajNhQmWLthbh58ME2wkKaBYx3
1jCkGYZWSpHRt1JeP3KQ1bCLf0YSHeOx1K2YFfoo33LTzMtJQqgQS3MH/RTek1z1eGV/FSpYg3Vw
S43TKCs1vKCvDRabN9Rixse36QcCuW+CH/uz+VVtpHW0FcHI9C61+FGHAUIB9iqEUiU08++4sGnz
KgPxY5QhmS1tzkPOkzD2qGjieJTU306hQ5MY0QvzWxmLswC+s+cwxeyTYev7TaDNdNyP5N9zceX0
g5AlGOeV6pwRU+lWDo88JMjdNquzYAKfBsGoj+LzTMzoPZFdiCv1EmOj0/yL8Ud0zEWx+mYVh9zP
xs0Z3MrjBzVrLNEw7LMII/7PKg4F5YHNvh1fM+3abipSav7O0OfYKzOUNvF1m294+Yvod9UT39Rl
+rkkMesgB98FI3R1LPe4QyfNfeVKyg1QkRHA41bzw4tZd/j0BjbvQ3Nc3XwCrGU0gJNk23JJtfVd
pn3YLaGU1RwmRqi+4pNCr5AlWeKA9ijTxphCF00A6Z1/r2PM/FiSRSe9Mkq4A2aQo6trsjdXchFI
k4pFlEhgrnm6uQPEMduQQEZjOPbL6veSjFmKcdicpmaf5SmKjjaK6qBOkpnSZU59HjPOYwCWOsV5
zTVFelLqMbEsNJWMF+jBHCJpMeyb3/RaUmQkBNvO1EYI73TyGLboihaC+qSMKuROr0PU0xK70RXl
RHFyquuinsxlbO74OCGbVN6vRiiSkHxrGq7BkOoPq3bV1r05F9/ojmQQ/UQgBL/O5d8nXyDRj/IJ
HJ5dRcxYciB03COhGtCmWIAuLOPlxFf6lB4Ui6+pe/TSjxziIlV7bnkXecVdo9MD1/5kOSPXZX3y
qout1G0OgKjtvpwqSt/w7ep7xnPLT+ePpPgsvloNuuZfJfavmwWeVON878Vmwd95/KwBtzTut0RB
acq+aAr+E04YgzfTagb59v+TI64YTUJ7EAWJkGKye5NFcemLQl+xyI0PxjhedTzP5aInoeo6LZNT
WBnTBnkvdqQc8kPem5he07s/xGxTEdMya9bcGHkNCbCF5xId7i34Iw5elZOuSA8sF9ji22r3g3gU
fpWYRGixORqCjzv5b6wv2BJFMuSDA4vZwc5GLtae5q8lajyA8h3HRA6USag/4ADkqMpPd57ibZH+
7klOKibkZpSKHqwSsMsmjV6i6M0KFZJWiv+32zPZMlNtJ1epDubHTFDBX1HtSbjlhXskS4xZmP6K
G4NujRMHaKevZHXDg6oyB9fB+XKoRcEoWScTDQYFQlMb1ltP8QJoeIy+5VMO9VDmaXOamWSqpOx8
QiSMzgi1zwmEaQLmh62yy/GrbbSfPe48Vr0iLH9lOInhmD+aRMfWLx+8cAyGwh8EqEn2eFhJlXP/
2NOf/w8e2btuYr5G6gYggDhps5kUGXuavJfkUALKVn5Zw5wFeE6o0EFZir5aA5EbG3/VulNPdA6/
iuLR0J2Ic+r1NU7lbMrWOHp/MDYFDvJT9rLkaeaMiGKVgsYrfHtqzwNhxCBwDdNMz77NDkwwk9Z2
cKHdOfTtMu3iZb58PzIalCXfmIPhi09PYCxH/zjA1M6rzs+jCiwweTTfQLxqSmG8sgd3k5GH9Isi
3O0mnSa8iCIKOaDWyNiyb8/MyBJbqtToQcGin+Bd/qgE45rCIXsQAbORDVRw0DxlBl15BsUMnzBD
kFBKqGNWqs2umLqO29YyISbD1ieRGgnV9OPsTyuw9KlmU92tWYbC/2YGexXul4O0CCMheFkK4KQF
KGmDMoNvLiOz13ZP7SDrShFeu6fR2g9uaXu4KS2GRWN79x4Yl3UZSlg0A49DMXAXrOhTSQTFRF5H
OL9N6TNHkBmf1YVxfz7jUQMhPRkg7MEdcjF/TxT9O9vsd8/cKM5DQ5AO9Vlx6lLdUqeNexWocsFJ
l+PcaXZ7dQ5wAn6cex5uDVwWY5qbN8r7NakX1shqb+ef1olEWyxyIfWMv3WiuipHeoRwFb+fAQJt
UOjWFTk9k9hRLR1KY+vgsN+ROvRSN1lYli16WCa6ELbypKP7UxoAUyXBO/UUkeYpu+yGWEqOHgyz
unpqLtSlW/LHv5WUuOyKY5bgE2C0uL/Jq7d/RzUVxdOef04AaVV21sS/cAf+b6rgNkmCvcZK5F1/
eg8CmyqisnEZLoKjOG7a8kckNyLy5rl0iI+epVOl5k/gT+w3gehoLYR72fEGn4UbKNOBt9G26n1p
M1R6aHoCb2wI3Kg4EEddXsMCaaNONxkOP7KvFvBRIKBiFIyHHDvLHxX7GhLrFzOuzQkbpzcjVEcu
JiYVJMjMFoUXtfNRfYIgfDFJdUTmx97MWzy3hbyaYnwhtT7zyMmZ4wvCGO2En4TV+J8Bdklh5Dx4
M3qPDANOWunUcckow10UYLI3ewq6mFAcOvcNjYaP3attk5WwCclqVu71ap2vHWSqqYtVh6b/zJtv
x7XaJAHMNyAnzMNLURVgDB+7oJDzZmY9Xn3xz2UewvDbVHfXiTiAQEIBYSLUXixpg/4oq1LJ1EYl
acIhSARV4x1N4+XmBvesy6BEzONr96Hg8tlnOHS4hNqGAhsT680yOuHax1dJZnybH2y4tTE11ZTV
0V0lvpiBx8EnvQw6rzqc8uB+7Xs1aFCQmM26dWLn5CHFXGPEDkDB8XvhdFG0HHnDzaEI5s97bSxg
d62oNphqxNizgSUiDP9gRsamOxS70GHL2smPMcA55fHGTCW5BxYAfR/XEx3fOjQjT7/sCjsIIW+h
2W5xDv5lkflXdvillYSlk/fhmjE/ZRFwA8gRoIWa8ysTTxZntvJl8LTJDUB5hcFclKKXLWd+5UWN
IkNs+V7T1VPCVEiyDFpF/3GwAbL+H1u0PYQVvdv4wEgsBBvQdbAAH9Etgt5hvCVE54ZtX1pWspsj
08shfS2bzPoODzxru9L4WgivQ+qFvRFzCxo12VFb3nRuY6EzesQ2sekJsTXGwdXe4AnANQ9uH06d
QvUmfvoS4HcUXys+nqyU6nw0DLD0bhUYbYxnQOsbzTNIoi/rYnP8NPh6gwKNgCOjXWz15lOARCoW
yzEifvzXr5kb/V0t64JXmyu4Tj5NimYWY7YAvgKlwcJhm0lDAi98PkqvBKhvHRhTUbr/WyyvU4Vm
KVN5CK61bmp5TmOn9zewFEmVyjb+z0ksWtMoH/3HwJ2MsgGCf6KKvd7UJqiMQWwZh+hraK/NtpGp
4ybsfU3/GyvA5UmsTnSQNoLGgntr7T49gfVX/+VZ/lrFtF8a8x/3FAEjqb8bpr2BrA00IE4ETGQF
TODwo54EVM38YuO1AuB3ZgXtQsHXdx733nWKptYgWQZc0PdCR08fryLAe5GuQJ14XxncyRoRBaHt
m5f6n3OATNZyDu/hn469BSLvdRZ3O8Plm4J44v3rlKBLaORtlXLHTs+WU+QyhMmnFdHBxJXEFlCx
9s7e7tZhnL33Mc8xr98Z/bFdZHJXIU9lEuiWWFXyzuOnyss6DntKaL9azMYfTSbv1VxLrnSzbVOs
Rz68rltvQAcWWwoU518tF970A5VMH7aqV/JOwiT4vR+YdKAHmCuq6GyY+7CryqVIrEWwSF9CgrYh
ObJO/rdDfZQRx+0BhPFV5j/NI53HyM+MSF6TTWpeAnUYTLdN6LFXrYdBZERRBkXWFNQr10+BwrKo
8tMubxMAEZHkA3H2WjPpUCxHcVZqu9FAJ6D7QLoi0aA6+q7+weJJq/MFP7F3iP/7J46jRyvgniXb
zBzkoJQLXWfJL/UHKH5QTCClPPIqGiymLS9uAI44657Gt6wr7POfxLgoDfTJ5uavfXJwFNh3p9Eh
XWRt+/+u7kwloqTgjogbOMmDtCDW6Q/Etwssm/MqHBLTZsRWHCle3JxoWhT5XMfVltFR0PCrUS90
Zm2OoMrYKvLiHoF4upb+37T1qHyI4hAetq1oMZp460/VSShUUl6TyIa1vzhWj0bFmnfEWqTUVtoj
RUf0Ox5KTubvbjHr9t8mZcU/SPdx8e9XyoOljs6IfKnfq7oBW8q5L/HXacIclxbQnliFA284exmZ
g2mSMGk2/A4W6S5MXj/QuiIdmcpuINISkr5dHHfzSwW6WB7C4IWIjdVhhiRFsahgReSyERA83wIk
uX36EDT4eE8mkn6Fw8rL7scYnazuGJhNjT4CyIQpzaCDae3NYBu+1LgDTY5zEOrov47Fe8fyfqAg
qwGlTY2MiSAAO/4luhj9dpOLRCMlv3S12/a4eElHYRFkPjo0kiscNGz9cT9mrRy9NaY7Bb7/SZ+g
Qg/xX1pJaSiFnCpth0YCCUNkh0GQQbdeiXbHzysyBTlSIiAp8a/7C8iji08cptvhpa/J/tGP7y+q
t5Wen6P9y4RiQjv5/miRBFybRTpm4MATl2l4Xzn95bb4BWa5B0Q730AosUBrKRf3GmV/L3o09/Ma
jHYHhZXZS/harxdl0jC5JD17u1ij6k9wDqQyn+niSXlBRevOPPz9a4Odil13LLZBv1cV1mkOHzk/
2386qa7vpD2PFnVClZZkmNUhUkqUSwY9PFMu/osYiCyzQrfpOh855UscwaD7Gjqw38tVTnddiGB7
PGWr6JEMjzuarazlUnina1gnOOZRq1ZU+Ez8nh2euwlBaHXE9juwRNEji5KTusVOentrYAUthzdO
pkKagiC0nJrjecfaDsHDcwFl6rVsirRIs0tYs2+jNW+nlEjr49JzbbLTA9RX0meM8VuY23XvGVzI
yB5gEjZDK7IoRbNaKl632bFU1pINm+AuI4+1iNZMrlVCkFiXeIDhGvt0segGDavkAebeXerEYUVG
WyPjK5Qz/RO5JAqCcrAxugqIVJViYsgRpFmgfNadDA5hBFtIWT+noUhYWBy0nKNHmAgk9HB+ODyK
5PTpDiGcIgM8kGWAIx16Bz23QOz9Zz4TUAOrnqKkyDynNE3E/9MtodeCdVopUkQq5zq8yh2+Vapg
gzzi+qnOCD3rsY0XMA7BZAc3jFa5oiLNItLiTN/q+NR9UHKihWXq3wcXM4KfdyTfmauzx0vbzj68
s5gbwRNYoWR3Nnyp63MIw/0nJMP7rchuqyTrZIpWrLsI7FRmUtOGhax9XSWiukpJ1YxI8Igj8i9q
V1rmjO+RQDFJtMEtf9ZJgF2q1o2ZJsjREX5YiHTlbPqTYDsBT8UMs4Jf+GfV+9QuqW0ck0ckyywL
eqH2yKeG5EF7UOVgk+9h4mgm1+bp4UuaMkKr8R2yrmY8rLWdZXdzYiexVz+FjbOoWcNc+y8U0zac
O9qDVZwedOrLYefIbkI+tfIbsAlrrfP4BxEeOOcfozRFL7WLV0448IExBcCMH1Wm9tMQ8q61b0+y
Vh/1oque7ptTiB6StQYrWOP48WQKJPiXubudUQkljiCb+2wHAEtiVE7NLPnSijh0BtFN0aoIyTis
Wp8vez9BDL0UC13KyYlOhuTbpAOpAH1/x6aiak+bi+mhJplIO400Duzu+4CXur1QmPjWiewT5NFZ
ik/gnUDQtFfAzxUfAnNlhnS+YwoMP7EAiT26vmKevztSe6gnFM71QQhk/Ls+mJSpx2BHOkwG/aJG
+aTMzh8GPORIfGbm+jQq0l8Y9N2XW72cZDGSAt8NmCWJBY0lwMgVntgVFwZHZs4ta8CDLGuDHBVU
rLg16lLrlGTw8WRpcuMSw8gQ/75zPbMRrXKEPkN0SH/N0NDb1sGMav5y6j4HYfexYLLvUc9dEZ6X
85qWDI1+bE8NyteV4QlBS7rjOj9uJ+UGs2v1HRRY3N/bVHYatvob6KC3qTu8jkw1Zo+CwDg61gm4
+ffZ0eVgdq8YKW+XNaLhEEZo3mBKsaafCmhY4qt8xFxsvRtvhPe653wDmNb0Wwa47eS8NYeKw8P5
EOooFKktKcW7eQaTDIGPJanxgoBn3s4tjlvmbfcL6yGdbx3miYVA8noT3c4hb+dnkflPTdIsVRKs
WHpsxZQlBjXeQ7Gn5Tns5uju7+Tq4CzfixfUHYQAWGReBpQoNHYdklVJMzuLILYBYG+ELX5eh3wG
zd3AfHuyqhGmfr6NTa3141CwXz33GS5H7eGwNWkJOIHtSgljwobx5xZpbCy34XmrhJPvZUQQrB5z
pw/1HbqlZe8CPK6ExZDWT0RISZQrC9GPzm/AJPbSuqcrgaQ+WQvOt//amhKTd651uEFeST1tV8ob
wq33IUCDePjC3yOnEs9pCuPydlEflz5MPItQFs2iz3zVXSo4ByNuvN4GSdInHrVsHrsUMuw/yUtA
slNXmjqUvjSqj7UFaKwpf7L98KeLd5mwpgir9AynHfsCnD4DLJCS3mg2uKjmwrxR76qmnoxZ5HR6
BSRu3nSNS0pzJZKxXMeKSJkdXMHbT668GDFoWrSUn0wnTvaGFUFzNfGqMH3GrYerfykpjqFTLD/T
9Ey80CBe/uuLYzV3kkNJ7Qa648dDMKmgZoGSuWwdKaWR2bDVy/MI83MK0u6g6LLe3T4wY9MfLnpS
L3SFN03T4xony0HF1xKoAS1agFxSr4eZsJgQWuU0+zj9TsH/036BYGirrwuTg+xtSu9qLSWlu/GV
/PjLcYjTdTYDcLhAa50jOZHtvjuTCRPgyqyzQiJCxYVLOegwDO2FQHKgxrRA0lOVyatcM9d5Wy+p
Yo+WPvgDQ+xtjSv/JL0z9U9dLulIzldLUBQjkWCtwtiUBWc2B3hJ+g0ecBBKL5ytoVFKuLi5dgCz
jeIR265lyHkafWc33oOptoeCZnSsqokae8/di8tuKYyOTDFQj7Ei5pokpIle8Zl3mChx8OB7DOtr
UYKpuO6e/gqv+Ij5THpQEhZKuXKNQZ/Rq83LAfB+8z23KIUyJ6w5Ej+flHu2dmTkFMLY+nuW/oAn
vOilhvMKxbZc+fkiGFk2BvqJJF1ty5/7cf9cjnZY+NxuY3dAGhSF6LzERVwixJ+eYwqv+KHQf23b
7gRz5YomrpPNke4Me28r+PMDWBMrvQxQXWS9OA+WOyGXgSExLTVEySOfVExcCy4b6e7Pb3jyxGLJ
CK5XK1X6PsgjzAxc61iQKboUw0/6CuGJ2e0BGI+Fwos2oge31k3ys5ZRlNQjJXbiKmiDCG1VCtnU
JNZ/InEYQ/WA6FDSCCekKK2+FLYssj3/L1H2wvKVmny555tSQXP7dPGGZtr9qvDaEU5QvFFEw1Ty
bjoiLOzrhaFSJ0VVYSfRAUfcEVO3sn4CRtbdNTa0BNj8AzUSgF+rLNSilKUlgxaLRL/I0hwPKqZm
d49WmyYC5ceJbGRJYTtY3mVOB8LCBarDQ5EiFElWgwn+QKI+sgsQc0OO5FY7uhkfLJzWeYxP+fjL
icqq9LlAQeGis/YdoOm5AwnZFEIF+d/zglRMdDowK5N5Jp2+U9z67P3yWJME6EOURrcBKKA5bikI
OK7qyhl6dT1/0Extvt9UHGUD2WqSMwB38KAvel1RP7+7FkMKKuBZXSltkgGwdwnOIKTHw3k4Z3Vt
GFU1yakkHS0OJQCsMnCxMGxNWVz8FF4fA28zXaIjymoZdbg3aaAE1xaY4h1/2YbTskBSMRqlH0ih
Jm5MbJS31GQ+78W9iDIvq5q1/d/GJh/d0JCYDauVuVSS8EAQFKAJWJ8G4Pz/YkdI+4nVX2MoZ/au
NbOJm/u+B072dfmhrLfsYlnHO7Kff/vZe/jqPBSs9wAo9chhewOEhNmBv+2xA3Lla+Pu0kp08EyG
iju0nDEVLwKR4zrXPUnS9uh93DszXIXIVWkQi2CCpzXrevAHaJAtOxCVVt9VjGxshTGesuiuaDKH
HKE1pxmL4Ls9JBOL6+8JwCrbQCPPcLY/qQ3PNFGt4zZFrk1rzAFdmJ/jTS6rRIhE/LQCIf1+bjel
xBug0nIUo9K+FZ1R8XvRU7AzmEiCz6T289+EMIR9DC0U17QrFHDFZpA4O9sBZ3NA8+a8NoqlfBFN
0rigF/hBIjWh1LucPzWTtXh0s69gMUhGdLBte7ciJmWeu7eQX3bteA6yaPsPN+BcktE/eEN72KLx
r1goVATqsK8YVjUJ7VDPfHOl2bOZi/fRpEZVxG1FP8mePghwsCgA+dJ4OOrkY2F8HTiMQ5q2FiMd
yvBAQlf3poBhKUkBdlYvDn3yqCTEiZJh09PDstGuqQ8zyrz4I36N5ufkONItHJBxzzpcv+RP1h1D
2EIMCPtKDDnJ5Sqa+/NelSyFG4KqsfqepUICmFjuQ9E7Y7Exk3vtcrY2CKA+2BzH7GVPMNwuKcfn
VXB/XDq3fkVvFXtfc7I1t1fjlAUjxb6wuDF6nCa8IaTC/qAHanTuCcbsqp+HTScUtWRGJEb7NGB5
i7CzWma8lPpz4Tn2/IHu/p7CXp5rNmQtPgsTZlpgsLzI/vtYxjJzeuv1K8ihDRPJDyhwIcdpex52
Pf1KoKPSnkY2IPGBQsv7hJYs6WERSj2rj+3aBnlDGvnryDPg4tcmkCZAm16RZPlsGhbiuEaxrXvT
ECIJgQy7qlcgNMXCY3OEfH6Itw/CC9fS21erLEhbVjt5WbikO7yf+BgGPMJpzRb2XLWFupPGa6hu
SBzjBy3U3pxjWiJAEAfXWejJqG/BSk6GVhZKPioLTKZ8G1Wz9lWLmbspsTRj5MXEtfnqkczXpx6h
/oMNc8cbJqjf7Q+kLNouBR0QKNx7tDAeUr/wk5J09X7Au16+K3JEaKR8a3zQCWpW6rh9u31kAp+A
rYhA81djWnrijruEEpvgFhoQGnPX6AeI6t1ZvVu6zVRDYcMztFwS/TuiBVlniRwW2PPwV3aY3gXY
K5Ggnlmw+cXw5IWv9i2L/Um3OLY7dVfaA3KKfE4JOWrvjEVdZD1UIj9adTk4M80xGrBky4Eojvj5
ROQ7XjDk5odChoDZSxOm/cVD26Mn09zLLkJmZRpA3HePyJZJ0DLXpQePdzCmoJXQepaWX6j/pMUz
L220h/QYIoECGakEECPXJAFsmNv8dg8hog3pfowRG90h4gWPRTXsSIXZQAaVmCEkki+9s01wWbgY
7V4BW0Bqtr9wtj6995s+JQWisyJiqtm7B1ZFbFcMqxnZGCN3ceSiHtOldsc8PwGCbhc4vs4C10l5
YhfDrmhY0SzMfsrM4mg5Hpa4Oh6ahRAFMUK+/ASiPajPr7fojBAriTuIY9kNwS1vVYjxbcD/4qS1
aENvUaSNb1crHUMx9H8QqyXWTR2MmeMU9z/U/W3l+6Xhc0nBaV50CryRBWqOI2Eo6wopFsbvvMcT
CsFWnGng3BFlX+3FPxDNKGRu47wfEt4R0Hr09PKpHCKXYzLYXwYn9jKHAWSvwtKsMz1MvA+MfVN6
XuKeheALQqewFHBku0d90bnodv5G3qf/WGycS/5nRaYkuORmiiqHSABuINrj4poCh4G8g61y+nRO
gwueDIbePPqOOfcf75Nkklspz6boJQKGMH4El8BMxFH6MwjklBIq0YGzC1EDNTaoNmX5io/OCgmz
QKBeXKKNNx/yZepkAfYr3oGGhXYaQgSS6QzBW1LkY4RP13YnwuJKIYuzRnYf0N+S9gE2dGkZNrFp
+M+xUjfUMLcQasWaIhpiogOZEG0LmEKILHRpizRWVrZ9UoZfwDUDpW2h+Efi5ILai3GK3fa4Scnl
gQmV32gUuXoIE6PtknJCCwJ87Qq6w9UJMBaYW2GRtdZxKEHJZ6IprwAm0r/uUgGjPU08+78r0KKW
CPOQsyPPepkJCIejIjqyJYLb4qrtBdo/7E4t08E/yEy7ubWuUis4uGxBGb9B7tvmgaHolkBkv3Hp
7dSkhCfbWrV33Vs76Jnj7Unni8FV82cghiTRxc17ZLnjMElExRxprw0qnF2EYYxaD+Jbz1m8Ogy7
r6ABrv/yDQWO6Q79I7c+1CgnwFHsWtkMWoL2fwQLxHNrMQ4pOWUnOBqQ71C/fFAx7ng0s0XqItJP
J1bHs2Posh3sayOJPxPhuUaUHjbeYVziYD3uu2f38Ep2BXQpSRKOG4550VZOMhnd05vPFWvVQAl3
9Q82KaE7GtdUaKg8PPn7UnRsfnGtGlA9O0Vj941BEjZNUJrs0oGGRROmNZ29WBDkpgiRY88zkvyV
TrajX3KlNh/LGwgTtu3CKcDrNfFnNZD7G4HZZcXHZJF6OGFW651v0TYEtBXpdYHxcx4lQ6x+nTGS
Ex+3spILifoNDOuEJscOleN0clHVYWVd73Jyp9oqBhrqDVW9MWHS+1mq1EVDE0/RvmV1OcRFVtXl
hJIXr3eAQiT/Ur0JTa5JNGC9sVyXYqfbzduLWa8FBUbEvm389tQ70oYZVr4s7U3jDNxD2uvujb8C
j9C2ptg5x7w/sgyGBzdhISyqOXQjl+OS/1v8sWLaU7YCIykue1PXFFMtPxew+TTkoqbsq294Gc6Y
cxFg496O7cOfW1h/IFfEe00qncaCHNYwGZEgwg0q1SsuuleMxlNCzfZXk2+P6f8eZJcsjOI1I4EH
2wpN3Zapo46Q/SR/lDKfaHpMBX4WzzSbsHBluduOU31DiPEyHFb0EO7fXB+yYdsAhE6A2/xWN8o6
5IdpbxO50hU1OP4x05sJPhyLcOV8M8YO8DgYcKJVpKWQ/4GuFp/uMsbPlDsZ2Uyv8NUEpwhVY2kq
9dZrl6pi25SLfpcGyJvB9ElZX2azWP3D4ApH4J7t4hU+V3It/opAhyUH3YKHJ3+vH9xyioqxr+uY
8XZGw53RISikR3gm+EtILYmRFgENKcStwJycq3GzNZ6Vz8G4IPLCDvNNWJQt7cq4PPVseSWlZTDK
qCISBOWUt/AUFLmIPXTB5oHEkJYrpVHcV7hbk5jb6WBrT5UdL3jz92mPJg3h3zN7Z02fQhdUim4C
YxDqj+SxpSt6WLoYKw7zhZzrC5i5kuIX2bIzg7PtjaXGsCwE8/7PRU5mecs4gDOre6A/GHAqvakk
M/k++WOJKE7dqNBoEJcPFLk3a3K3qXiFODK9+wjN010ZaCanMKriQRby9lnZCdzg9SZRGoHbjMNL
zEhxXeKkUI8WDxOZaTR9gL+mCaoGS0tpNBAYs1nfvF8/BsHnr/8+oQuWbTVxo992H+z6a7h7cObg
E3kc1MsZC7tYzQ3+1/2iaYcLK/xWWHBQcjQQ7eojR5f0JHQHMUmaawv37KvKry7AwYDqhe+T5ucj
btVGVSRlNZ8cFO0HndB47BcEk1xMDw7KJpj4y4F1dbhqPIFSHjOgLJRnCDTVuohltm0BqBA22vZt
J9/ae7JGFt0QbmLsqsWOpv5qavZQO+OJckS8f0ozYFyzy75bmrGENevPe+FY8Skq3gX2mhRPIKnd
rIYBhbkH/qnbFdrZzF+a2Yl9eFVEIydVutfA9JK4l7fX/kYFhPCitgmACgYO10YdRf+mxr93W6Ej
YZlOASRc42kNdsdzPbdmyFE9EfSPIUKAt+29n+KWcYrHHkhEr6toHk114ZqTMFZZcqJpaVwoi6lq
MiYRAT11AH5mUhYn8RqYj/aueITShgr0JyXCS+tlYNNEWkfo8nvVfcDgyAHuGSC+fXIFvpZW2PH7
VINQrIyJl9J354iodcCInQr6nNTQV70NzRnmcyNe1qyHaLmfH4uU8QrJsPGoXcNhL0PS9M7qioGy
8BTZDq+4LYjmB78vuuxUNkynU70OX67/h9IQGLLidXmPmzpNBSFmiq6yd8uaysxoTwSH7qJEl80U
RM0RpzgCz5tt5/hH8CrDRk5cCItpi3Hs04m13G/yry7Kz/e2OgKnqHF1eP0UkU7KfeLLtV3ie0Nk
uZt9/QmnVlfWMIB9lSTHi1atKix/d18Am8aMVhmQFrYbujuTDyuQnDj1JJ8iQFVUnd0QQaAi0TsJ
Lai577S/iDvwKUS99D/L+r44J8k3y98Sukc9pUSmQn/b1itc3JGPhWFo3WbVCQn+hmsTqOy5AvCI
XU9OhpG759F6grdjyVwWnEmFfSUATv1xuTpck6cq/yIZAtYDeopT64kYMztsB4IoDElBKZY3/gP6
z094SsFtGdVtiXzbWawRKOgjUgVpH+RcLO7Hj6PpILfoZumdnvWjWRkKcYHvDsmqdwtkbIo8yJCG
OdiTysD8GpWcgthGf+neJzDf7VfoHwfhMxPQfIT5DBJxrR705G8/aLYy0HJ9ZKSE7w1KwQyKrstp
HOGuexZyQ/ejH58UKoses+nKiORgJILn1gS3xpE1tCFzZFEIhLMJHRtJT+gOk/mt4/qN7fDVx5Gg
QMfegm5vXLFMgRCP4NAwRpBGUlImrlUIjadUH8Wvit6G1jd645o6iJGidwx0Tr7/kpiPd6yV04gB
M3Mx7I/Yd0KpGVue35pyto9E8iQ85RbpAwBpuz0Ee3LV8iIJBZci2GjzMudLQXkdsnkRaEY1J8AS
fnT2/DjTVeosEPm9osnp52jhaqXYDSMHC9SOBRHfqJQlR0ikoCrlgv8tPDD1I3//AWyLdNpkkvpM
I3ZtJdPGq4bNigWRnaN3RNABEGSFrPlOeDb4wyUvjbxbjCpABBxaN1SoZnQoLgP7n4tR9ERcczHQ
pJdWTHdAn9ENjOfF8YYyGW7itoCz3O1X+02YYZXhkzHdGBESWcnHuQfBHSeDYM23r8JbwOrI2N93
4SGdSW7H54u7YytfpnxTbVvfCHdJ4wkR3QaS7JAENicmXotxER8G0qx9+AwQMmch7j9nGIgpqUHI
mllw6AUcXDBZlR+iQKI4/t9fwK/Q7V3ZrPVjG+8s/CKEYqI+LB5RkTw/s+ETRKkhYmr8Y0e699Ej
TXq2PsgzhuRQg81R79d/BokYIXFF7DgPy6uspVLzTMBq4llVZRZk/eRrKKRdWLzSFoEApPQwFtwI
NrHPWo2w1YxqUzxogTHf+T7RKY/sVY7jRac88o1WMaT3a1Wxjme0ACm7paWhlU3dF1Pm+1074Gpa
62pmq/yaXn3tvK+xy7qfg2F0Tj/4EknYHmndEQWO6hnxeVdLmFV7niGpILnlcO5Wb7eDeA5YdN3p
ElBzCNxojH3/gANq4L31vHMJ+K3B5dLSJ/nGSyFm4UvWw1c+ZIOFV0vEXFyZXAhmZg9CuR2CGfG6
AFrQeAZAUvubwThFYVsLeDollJ9CITVRRW8lO447Wn9XtxDiRCiCSAKWMjUEUPypewofFYRee8mG
N6OBB3QPrfVv+n0isVeXG0w0GbWEVFoB4i4pswjwnDYGdACNv3Xm3c0p6aKV6R10/rTzWejljXK4
cAgEcgByMhbeqeVj+PZK6HJCmTGEZjn56veq5/EN5WYvsrmljcw5zCn/MpEgwPXaWA3dAn/GkaU/
3sNQeWzHrt6c2bGmhUiTaLpzXqYARvRxzkK5QA2uKfc/LUZO78lG1weucGEKYiV8c0grqc+EJLai
TsAAE8bRAsAIDHM9rBhOVo0qR/+bcCtzvhLfHCOtuSiZQ4j9UmMyM8CC4Hz+xxka4bX99XpCbElz
NgpyAjmOWENb+sganloTYaPySkzO+2faiwoEJIPmhFX03pwfvlyYRkQ9/huAw72FaySIRGWF4W9S
b+0FOidEg8WMg+nbgDXz6CzosrgqI2S/feyvqwhX+jueJ9RxSGCPFgmQCVuEMpoaCAe046Nq20Ua
aDoJIrv4+n93dlwk2ahqbzhvf9cMmvra5jLTueC/ianOzhmi6EJhch9IsU/QTa5xPmEz0YhYfq6A
L5O8Hr4r14KTB1TPK7iAMc96C36zuHdE/5WdQ9qACXgPTKEDYC9zCrm67t8Tu83r9/xpveuJ46eF
QxyYeRUrPtQ0Ci00Ea6IMmdUz91DRXk1U8gwFD/wBlhiL3iPdXGXnEKxuGUBEm4mdPV3R05eNVjr
m1tn9yncVj3GrCagwLw67eeqZeVGDcmAs6jxCQF5qaa80zQDRpYEcMUmSItT93cdcEQYlOkvtJG2
11ginq1/H6/O6DpoI4+DX+TD1+XQmvC3uX9FfEEk18NTEyImf/fVHDlaaFj5DXVh78E3TX0t9hDe
R/q/+wEN4Gxl/995E1ctiElURRscBOc1d3MSK8LXG98YhEBFiFyarEX5JjXd4HUj5lofn8VJnEVQ
yWUvx0m1woyYXsf1MFYBqwwek5HSHL/qr+bYHmDyuA4BNeCT5MZ50ZxzrvxwZ8ihVGEH19feyRRT
qHTIN01TR51sFX11xwhgGv8fuc7cT7BW1+Dt2cf+UGbSkhgZIg3oT2RG0uDw+yxB1/lfBCkk08FG
w9lj+repEKqZ9s/SFGkSxSrvPkZG4v5nPdkJ+USXEpQKTnY6H6Ev5fkO/w+T02TEjuj+m38HXXFC
eIqvsIAI6Bp+Jnm2wYC+9fwpSjlE8BrTXVh6kGPp80ZdIcYFc2vY06G+DGBQZfQKy66c0M/AtpX5
nGwinGk3bP4fPTH+gwvsgiXsqI5PIOIuFKm0nAELgr3Sjcckv9PO6qhFS9nwAR53Njlb8fGYyE+F
ZiAjCz+6ojDYI2Az4+KNBAkr34bDPMFQ9UAmIpOn6+aFqDMokJv959iEbbfbJUbyByTH4MW09tkT
jr+TiZZDuu47IL91G+r9Skojgb5WQLdGaoWAGz51dYPFKGRbsr/siFXgMD1IXHVeaQ1d74zk/DGo
h13z8lwZiBvw8DE93gKPQcE8kfBnJWYQbuXkgq5BzWfT61xcGve28JZTdCR2eeu3FojA6aNxxtdC
KUMSBoeRoX1Mp+NjyJM7GN+lpYJNblm256hPeeKDOc6ZNZKkR0fZtxbXW3LYFufCL89IdbXymMDC
mQzNVw4hAviRYTDj/aRs4zipv7TttoeRmdwRHJprmmHMPYSO2MSaNP0Jd6k0YsWhMexqmYqJmNW/
mD1aQwPBbEgOWYgC/JUCz9SSRvS8+5QL/q09nEaP7BKRq0uMtVXqw69xQVIIZMyDMaZKnrCrT22l
k7nOLLDhnVQ+Bjmk2m15d3uH35hPnGmwvyQvcq3sB0BringXUDESll/NJdSvBjRWqIXdmyMELQHn
U7zodn4siJ+YD7/XKQBlQgZTv/Rhz39NZTF7Sav8ooo2jYUkU0cXgFzKjNA/a2cv3x7BtFrwowN9
rlmikt4ovJytTGGKTaWpPePONslZ7PeMy3P9ZuzdDaJvxBEKYFbqW10qXfqspmdzlLAHdl6doTPA
ftu9XrIPmUA22iJWECwfDEkeLyScPcnBML8ngHxICbsYjFacSI2p2KEAQaan7IZ0Z8bZ36QfcSiV
EmQ9qGxgfS9eq43P7pXG/THTGuViYngSNzUPcXW/LkO65Fja+D5HtkFBo0p5GRFpX/2ssLW2nfO+
bS+sX0+0MHqrTRDZlOHnn9+xVz3Igyb/csUCMljvLHwfB151A3Oi7AYpG6LWvign9kGYgnrbURPP
voikvTl+rso7sY0lCG5D9cAFFF/5UyORiDSvr7YvDF7VT/VxfaU2CfZA7JSQZqYf7VZPQQHvMZO2
seD0yUkvb3gsS24wP6YadsZciyLLpb8KGc1CedxYQr3gQeDYTXMBdK9HkVlnHJ6idKoRdr7pTJcy
twS55dS+4XJMwpqqQSF/x5ucvqodxYJP3TMxDlBZGgTgaBGq20e45PxRcnWR5juOjyBlNZTZlUr7
8Veqn64+VaF0ceUgmIleXPLZfkZdCvmvKgCHLRSS9+savxFEx+DXx3opVdpRyYpKk6Vu8demJmdN
CadMtyRIqqHOsGJxq7zh1GMiagkIMKn3Wgvh0x23PuxM0/RLX0eQyY08BaPvja37yxINhIL64Ae2
NI2/A1oicddY0oEQqeRV90A41gKDVhOHQpKHicwaW3p2q+xdHkxyA/UyyHOQ1YMmHbaH4vAymM95
Se7yeqVgMJ+KcpbsnnDFLIUTkeBOZXTG119NSlSlt/ra+9jDZhEmsjovOBTgr1CsK5CVhThGtXzd
JjAu2FWhO0NNjpzIht6zH7quuPpGXOtyRt/5C2wm6XTB5v3BaIKUqaLzcUWA9ymwNMuW/8Iugpoj
fd4NgjDf/gWsMyHZhl3K36/hr+K0enfpgc4T8qyJHVk0r/VIYsvNpc8k9Pgq164W60eLWKPVp0sp
GpQxeZJ7PAtSrSYZfb7EPXRGesSEJBzf+WrWzSIWuhNZmISm4AL23ysDQMgPjojoxdyOPRUaCIcI
ROAwWYr7wgGwKZNpRUBbTb+3uGltCcL3OPiXCtvAscwNRI9urinQC62vThdBe9BPrIui9DoJB6Tr
tzRB6gpUOj3fXzphjvqlp8NjuUBOXP/YERcTcTC85p+CC3V0ONkMpJR1igDnt7XDxYG1p3ojA7cN
6yyKUtn51rBzp3OV6ED4cAWDTg456JATtuTGWoAoSDscTBDrM95ceAA0oTTv56n4eOFCa49cwKQc
gUuA3YiDJ8A70mthQTUiSSL+dTtK1J4xWLFQQO7jSDqL7nStRg9tJghqgKqXQcItpVH94icpPrAB
qOg+MhnD3dmEYenmlDDYkQVdI8zhXne5fKW+sjkHBBTVXMZddQtKN9yUNAAAztAfOnIihlF8DMHw
45BftkDsTWqpb040f/SMf3qk5Id91I8SzFlOScOtcw+JwKfbdJVQ1T8/oVGfRw6zlQEq5+vpcMVi
kbBKtzB0Lo2vEyFQ1RdoBpmibiw3U/Oy1SVJyz9/6K8ZGwuG/6aqL9C2rQD7V4yGoUhagUMD+Wdp
vurMaWgx3vKDxZh9B+PW/5EM9xqZDAQpG4cZSjYG6X2FFXfbezTA6JT9cvvdsKlewV/svogONMbD
llZIFGYKUlKXTDHFfa+DPPU8lc9grzErf4Gtn44x8cO5OYGCEX2dDWiEZ9vgrNiu8PJ3PftjupAp
kMawNtFiJveQFbVnQDVQKQJkV68hUy/t4c6dpjUKCbrVJVSiR9tTt7gYS2iyWlg0HZAqlxLyi5qi
uZQMs1K4luZDbkzGdI8z0sTCV7uTv6MwDUYATrigg6GugDnFC++KlHNSioovN6OLjO6arLkzusec
qWDlLAfPafkZY3R5jGZlJCe8FYA11SZoxOoaerPgdWEsm5TxoiGfJVkZ05pIpvOnocU6TnIB/hLg
waNnvfNQZQHkg4OddZo35c+6t5q076R2RzV22AcRWM5o3zCRMQewuBQiP8/U9i0kCGeguthF1XEe
z8nsIlYmHMrqI6qgUVafey3TWQbQVM2CKe64ZuTR13cqo/y2zfM5Ugw2xswT1v+pu+zdH24IxX52
Ewi+Y6x9VpjspyNpbGBmgd1DhlL3g5/GTz3K50YoHR2WUkZX5jnxI5VZap7dBv+uXu4Yq1Bk8kWL
Mg1W8RB61uGAfxAL8ByhfCkamtjzWIJGtaJ10WMWKCAMT9B2H3dnWOHT4kyqsvNshxn29q61p01P
AgRsrunSK66JGB+KJJmppHUgWwFowSBu4aLK7gF53IR0bqnrNpwXjrMUmAUz6M5YpYm16rAb3mFd
/sRVjeGS+niPEeITg68PUiTQd1X2CdWg9+sO6LwotHVUaHuzFdR6jt9FPLChYGGBmm66kVJRxNvN
sGQl8Z+rCXutKJLoATbhbcAzvwG7FET6nFSfSSO4biMw3ltnVvM6B75RdY8Qm78EP0aYuFpHRbcR
CwKxi/RFrSHawhOh568EhT++W9aC7A0O4Aw6qvLCJ2NBBCgFE7RSokDaGSk/6puATsAdDcn1Wlo/
8rTAj6NaPzTVvq1Uey7KEMsuViQSolnHXZZxdAquuBSF6LUsUYrmNJ33CWtrDuTdG3qI6IUm1eXj
phOEANibNm9ERaJ/TdkrEUC5/XEqtSydLH1bJE1gF6/j3+Qcq383m79T5lABKZ/lHs5do7Dkl7z7
VXCiZzIyS00jXKZqj01wgPzlxaf06q/4hp6SmtGg7FnF6nAlJXk+YiTxnI5xWPveJAQTab1+3y4f
WxAqweKRCLulfS9E6cZ5wbfyBAx324MWMcD5EUZZr/sWXHQbERIC8XWV7+mMwibtrxFDRzuGdXGX
11L400n+cNSDM9WZDpKSxo4/YrL5IUD9Do7U95oEROKt+hrfresrVHpPMSM81qlk2x8MR0DAFogY
gaIUlXEpJult89jNL9zRslw7TPnAw+ZJrPE4vmdxRJgij90VS2vhMi/3NdzD0eIBLcrN5q2QrGKE
J/X5WG9jO59f9eG3L2uqKOPlAqrxtpVNYd/Ckw1756Qib/yEMTvj0Zz4BwM7tZvB2UYhRKgG0Peq
sW9uc9VyFK6lmKxNY+q0FxKjj5ravlBAZAIPOtEmVgS8QlU7tD3+kVBH+IsK77xo0WIJvdm7Ptsf
PI4rdBOG4NmSLhlZ4az1qOZYJaiJ7BaDs5Q1qzDuQGxvtbc+D1iWQ6iGRlglCqiEZmFirqsluAct
V5e5KoyhHmMMKmG//WjUB2Zw7cXD+AIjbyCBDug0ULD2c1/x7taih9+VOz30SBKzRpoyJubXMGlc
/+GunZ/c3YygiKKDPlo4zd6Nk//ZUD82+/tmsyBq8ZxCOz+FV4UbO5GdFB0=
`protect end_protected
